�s�Xo    �0 0 ���@����@@@@@@@@@@@@@@@@@@@@@@@@  @          �                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �8����O�V+                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo    @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo    `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo     ������������K�@@@@@@@@@@@@@@@@@@@@�                                  �      @ @                                                                �a�@������@����������@@@            ����  �s�TU�   �                                                   gJ�  �j�� �                                                                                                                                                                                                                                                   	��4�e_ǚ���                                                                                                                                  0   0 gJ�                                                                                                                                                                                                                                                                                                                                                                                      
�s�X ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo       �� gJ�         gJ�  � ���������K�@@@@@@@@@@@@@@@@@@@@�        ��s�`� "�Ф�                   gJ�         �s�h��                           �   �                                �                                      �                                                                                                                                                                                                                                                                                 g\>���\�
��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo   `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo     C�������@@@@@@@@@@@@@@@@@@@@@@@�s�dG         !@@�������  \������@@@   �   \������@@@                      ��������@@@@@@@@@@@@@@@@@@@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@      �       	I  	                                                                     ��������@@@@@@@@@@@@@@@@@@@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@      �       {                                                                       ��������@@@@@@@@@@@@@@@@@@@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@      	P       �                     ��Y���w�<�&                                                     ����@@@@@@@@@@@@@@@@@@@@@@@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@    �  �  0  @                                                                       �������@@@@@@@@@@@@@@@@@@@@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@              2                                                                                                                                                                                                                                       �����q��'X                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo   �                                                                                                                                                                                                                                                                                                                                             2@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@   �@@@@@@@@@@@@@@@@@@@@@�@@@@@@@@������@�������������������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@        ��c!��ݸ"̓                           @@                 �������@@@��������           
��������@@@\����@@@@@@P����@@@@@@@@@@@@@@@@@P����@@@@@@  ��������@@@\����@@@@@@��������@@@����@@@@@@@��������@@@  ��������@@@\����@@@@@@��������@@@\����@@@@@@������@@@@@����@@@@@@@������@@@@@����@@@@@@@������@@@@@����@@@@@@@��������@@@����@@@@@@@   ����@@@@@@@@@@@@@@@@           2@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@   �@@@@@@@@@@@@@@@@@@@@@�@@@@@@@@������@�������������������������@@@@@@@@@@@@@   Iw̌���V��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                                @@                 �������@@@��������           J ������@@@@@����@@@@@@@������@@@@@����@@@@@@@��������@@@����@@@@@@@   �����@@@@@@@@@@@@@@@           2@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@   �@@@@@@@@@@@@@@@@@@@@@�@@@@@@@@������@�������������������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                                @@                 �������@@@��������           
�������@@@@\����@   V���E��鬣�h@@@@@��������@@@\����@@@@@@��������@@@\����@@@@@@��������@@@�������@@@@��������@@@ ���������@�������������   ��������@@@����@@@@@@@������@@@@@����@@@@@@@������@@@@@����@@@@@@@��������@@@����@@@@@@@������@@@@@����@@@@@@@��������@@@����@@@@@@@   �����@@@@@@@@@@@@@@@                                j5       p          �   �  P  	��   \�������@@   �                          �            \����@@@@@ b                                                                              �� @      �Tm}�F�/%��             	      \����@@@@@\����@@@@@                                                                                                                                                                                                                                                                                               �@@@@@@@@@@@@@@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@�������������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                                @@                 �������@@@��   !jE���@bN��K�������               ����@@@@@@�@@@                     �@@@@@@@@@@@@@@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@��������������������������������������@@@@�������@@@�������@@@@@@@@@@@@@@@@@@                                @@                 �������@@@��������                                                                                                                                                                                                                                                                           "��J����m]�)                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   #�s�Xo   `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    $�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    %�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    &�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    '�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (�s�Xo     ������������@@@@@@@@@@@@@@@@@@@@@@   p                                g   6 @ @                                                               �a�@������@����������@@@            ���� �s�TU�   �  h     `                                        ?�G7�  �~�Z) �                                                �~�Z) �                                                                                                                                                                                           )��~�����                                                                                                                                  �   � ���     @   @ 0�}��     �   � be<           ?�G7�     �   � ��           '*,	�           "                                                                                                                                                                                                                                                                                   *�<��|d�~,��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   +�s�Xo   `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ,�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    -�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    .�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    /�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    0�s�Xo       P � ���   0     ?�G7�  � ��������@@@@@@@@@@@@@@@@@@@@@@�      ` @6 �s��U�� .�M��           
~6O   ���       �s��b��                           �   �                               �                                       �              �ǁ ���        �                                                                                                                       ���� 0                                                                                                         1��`4��#ho��                                                                                                                                   /ǉ������@Ö���������@����@`@����������|�����K��                   p��� �       ����                                                            ��� @        ��� ����                  ��� ���� ���� �                                ��� 0                                                   �   X   `  `   �  0     �  P  @   �   �                 22~\	e���-M        ��� �����G���=��'L�        ��� �������@@@@@@@@@@        ���  D�����9{���.�        ��� p��������@@@@@@@@ P@�         ������@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@ P@�         ������@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@ P@�         ������@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@ P@�         ��������@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@��� �      �                                                 3�*'}�o^ڦZ�                                        ��� �                                   p                   X         u`     `  \          u�     ��  x         |�     �`   �         }`                   %m��m���      $                      3                                                                                                                                                                                                                                                                       4�~<��y ݛ�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   5�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    6�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    7�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    8�s�Xo         ����  ��� ���� �        ��� ���� 0���   ��� 0��� ���� W`  � �                 ��� ���� ����                         ��r                                        ���  ��� P��� �@��� �P��� ��                     �                                                                                                                                                                                                                                                   9����T&ŭm�; `0000    00@`    �� 
 
����                                                                                                                                         �           ���                                          0�}��                                          be<                                                                                                                                                                                                                             :L�HX��1Ƒ�HH                                                                                                                                                                                                ���                                                                                       h       �                                    �       �       �       �               �       �       �       �       �       �       �   0�}��      �       �       �       �       �       �       �   0�}��      �       �      ;�qdD�D�R�    �       �       �       �               �   ��� �         �   ��� �         �   ��� �         �   ��� �             ��� �         
    ��� �         �   ��� �         :�   ��� �         "�                   ��� ������|�� (�!��`]  �A  < T� �!�3�@| �AڀSA݁�� @`~  �| �\ �<  � (�������_���?��c�  K��`x  )  A�  �} (;_���=  cC  )�cb  N�!;   ����^ �_�ă?��;y {{  ���)� A� ���ă_��~�@A� P�?���~ }9�@@� � �8H  {:$�*���;;��{9  {:&�;��   <:�ӐP4��ɬ�$;��؈�X �Y AՀ#K������;x��{{  {z&�;?����Ȉ;`  �x  �x AՀ#K��`;_��;?���� �� "�� �� 2�� /�� B�� ?�� R�� O�� b�� _�� r�� o�� ��� �� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���cC  c�  H  ��a  ����= 8:���:����] 0�`�z�' ꀁx(5 	|�z��ct  b�  �� 28�  c  b�  I�c"  N�!A݁�Aڀc8!`� (|���N� !        ������� u`        �����������|�� (�!�A`]  �A  < D� �� `�a h3� | �A݀� @`~  ;� ;@@@SZ�{Z ;  )��[  �[ 	�[ 	B ���[ �[ ;?�d;@@@SZ��Y  ;�P;@@@SZ�{Z �[  �[ ;  �   =������+=n�?�;_�H;`@@�z  S{��z �< 0�?�n;� ;@@@SZ�{Z �[  �[ ;?�@;@@@�Y  SZ��Y ;�;@@@SZ�{Z �[  �[ ;?��;@@@SZ�{Z ;` i��Y  �Y 	�Y 	B ���Y ;�;@@@�[  SZ��[ �[ ;   �?�p;_�`;`@@S{��z  ;?� ;`@@S{�{{ ;@ I��y  �y 	�y 	B ���y �y ;_�\;`@@S{��z  ;?�h;`@@S{��y  ;_�t;`@@S{��z  ;?��;`@@S{�{{ �y  �y ;_��;`@@S{�{{ ;  )��z  �z 	�z 	B ���z ;?�l;`@@�y  ;_�p;`@@S{�{{ ;  )��z  �z 	�z 	B ���z ;?��;`@@S{�{{ ;@ I��y  �y 	�y 	B ���y �y �y ;_�0;`@@S{�{{ �z  �z ;?���`�{:' � �x(: 	|�   >��ba��W/�n{�cv  c7  ����;@  �_���_��� 8�| @�� B��Ț������:�� ;V
�ڰ�c[  :�  ��  �� ;   ������ H�| P�� X�\ `�_�������������;��;@  �X  �X �X �X :����`�z�' �@�x(7 	|�{[�ct  b�  ���;   ����:����@�z�' �`�x(6 	|�{z�cT  b�  ����;   ��@��H:� ����`;` ��a:� ���c;@  �_�o:� ��p:�  ���;� :�m���b�  :�  ��  ;_� :�q�Јb�  ;   �  � � � �`�{7' ���x(7 	|�z��ct  c5  �����] H�� z��;x����� �� ����{7' � �x(7 	|�{�b�  c5  ���;a p��:�� �� ;  �  � cc  8� �8�  D  �:�  ���    ?�ǘNn�уe�*���ꠁ{4' ���x(4 	|�z��b�  c7  �����/| �c4  c  {�@� cc  b�  K�c`t  ���z��ꠁz�' � �xz��(9 	|�{�b�  b�  ������z���� ��� ��������; �eʪ{&�~�&t���� z��-4  {u�;�@� :� ٨��� ������?| �b�  b�  z��@� c  cD  K�c`z  � �{W����{[' ꠁxz��(; 	|�z��c6  cW  ����:�� �_��{x�ꠁz�' ���x(9 	|�z��b�  b�  �X rH  h`   ���m)�  A� T�= X:���:��m� P�`�z�' � �x(: 	|�{�cr  b�  �W "�_�_�W B8�  b�  ~��c"  N�!H P|�� �; hꀁ(|�b�  c  �_���} �;[ ����(|�b�  cU  ����`      @j��w}7n�B���= �:� �� �(|�c  b�  �_��} �;[ ����(|�b�  cU  ����;?�l:�@@c8  ��  :| 2�S  �Y  `   �} �;[ ����(|�b�  cU  ����� �; ��`�(|�bz  c  �_��:_� ; @@S9�{9 :� ~���2  �2 	�2 	B ���2 �2 �2 :�� �^ 6zt���  � �t �T �U ��  � �u :��P; @@S9�{9 b�  :` ~i��2  �2 	�2 	B ���2 �2 �2 :� 3�T  �W  :�� ;�P;` F{u��:`  A� 4~���6  �X  ~9�@@� DB@ �6 	�X 	~9�@A��@� ,:` {taN   A� ~��6��~X��:s ~9�@A��;@ A� ;@  
  {W Јb� �얋�) �@��� �:T �� �(|�c  bW  ����= �:y�@�(|�cT  bu     A�侬����K�����;� :_� ;%ؐ���  �� �� ��  ;?�0:� ;S4ژ��  �� �� ��  :_�@:�� :�Cװ��r  �� �w  �� ������z�����v �zt "�� �:��i~��-�  z��~��@� :� Ԩ�:� ���  ���z��:� ~��:�(����  ��  � 	�� 	B ���� �� �� �� �����������:� p��:� �v :� ��  �� b�  8�8�  D  ��  �x �{ ��  �  �� �� ��  �  �w �  �r H X`   � �;t��@�(|��_��� �:��� �(|�c6  b�  ����;� :`@@Rs�zs c  �r  �r �^ 6{t��  �4 �8 ��  `   �� �:���`�(|�bz  b�  �_��] �:�� �(|�c6  b�  ����:��0   Ba�gΛ֦����z; @@S�{ b�  �  � �^ 6{r�:� 
Ԑ��4  �� �� �5  `   �� �; �`�(|�bz  c  �_��] �:�8���(|�b�  b�  ���:��@:�@@��  Rր�� �^ 6z{�;[ �؈��  �� ��  �� `   `   �= �;P���(|�b�  c  �_��} �;[hꀁ(|�b�  cW  �������<��?�����^ Fzx��x  {{ cz  ꀁHkw ~��| HV �y�zz�!y��z�,����] H�� z��;7pؘ��X �A":��� �z�' ���x(5 	|�z��c6  b�  ���:_�H�`�zX' �`�x(8 	|�{s�bt  bU  ���;_�� �{W' ���x(7 	|�z��c2  cS  �_�"; p��;� :��:�� �x �� �� :� ��  �� c  8� 8�     C�S����R�bKD  �`   �� �;V�� �(|�c2  cS  �_��} �:��ꀁ(|���������ȓ������ H� {:�:z7`�Ј�S �A2:_�ꠁzT' ���x(4 	|�z��b�  bY  ��:���`�z�' �@�x(; 	|�{S�bt  b�  ���:��H�@�z�' � �x(9 	|�{�bZ  b�  �_�":� p��:� :��:�� �v �� �� ;  �6  �6 b�  8�08�  D  �옢��{�b�  K�|r��;�d�[  `   �] �:z�ꠁ(|�b�  by  ��� �:�����(|�b�  b�  �_��:_�h:` �r  `   � �;5 � �(|���� �:����(|�b�  b�  �_��:� :@@@RR�zR bu  ;  )��U  �U 	�U 	B ���U �U ; `�  ��  `   �� �   D�0 D<h��o`:�0�`�(|�cx  b�  ���] �:ZHꠁ(|�b�  bW  ����:����_��z{�� �z�' �@�x(8 	|�{Y�c6  b�  �� :��h�_��zx��@�z�' � �x(4 	|�{:�cV  b�  �� �_��{r�� ?� 2�_��zt��� /�� b:��d�_��{y�� �z�' �`�x(2 	|�zx�c  b�  �� r:�� �_��{r��`�z�' � �x(5 	|�{�bv  b�  �� ��= H�Y {u�;pب��X �AB:�`���z�' �@�x(6 	|�{W�b�  b�  ��;��ꠁ{s' �@�x(3 	|�zU�b�  cw  ���;A p��:����@;?� �� �: ;  �  � cC  8�@8�  D  ��_���AR����z���[ zu�����z���X z{�����z���� &z���_��zv��V 6zw�   E�SB��X�UHp��_��zv��V Fzr����z6�� Vz3����z6�� fz0�����y���� vy������y���� �������z/����z/' ꀁxyֳ(/ 	|�z��b�  b/  ���ꀁz����z' ���xzԣ(/ 	|�yԣb�  b  ���"� �zv�� �zt' ���xz�(4 	|�y�b.  bo  ���2���zP�ꀁzS' � �xz��(3 	|�z6�b�  bO  ���B� �z���`�z�' �@�xzp�(1 	|�zP�b  b�  ���R���{��`�{' �@�xzv�(1 	|�zV�b�  c  ���b���{p�ꀁ{s' � �xz��(3 	|�z7�b�  co  ���r�@�z�����z�' ꀁxzғ(0 	|�z��bP  b�  ��:�;�p:��`9��P9��@;�0:�� �z �z �� ��  �� (   F@߰��i���y��� 0�� 8�@�� @�: H:� 	��  �� cC  8�P8�  D  �`   �] �:2p� �(|����} �;s����(|�b�  co  ����;�:�@@��  Rր�� �� :�� ;4 ٠���  �Y �Y ��  �X �X `   �= �:��`�(|�bz  b  �_��� �9�����(|�����:�� :�@@R��z� ;  )���  �� 	�� 	B ���� �� �� :��:_� �  �5 � �  �2 � :�P;`@@S{�{{ bz  :� ~���z  �z 	�z 	B ���z �z �z 9� 4��  ��  ;?� :��P:� Fz���;   A� 4~���9  �  ~1�@@� DB@ �9 	� 	~1�@A��@� ,;  z�aN   A� ~I�~9��~��; ~1�@A��:� @� :�  
  z� ��cz �_얉��) �   G�iG#>މJ��@� `   �� �:n�ꠁ(|�b�  bq  ���� �:V�ꀁ(|�b�  bY  ���:���;`@@S{�{{ b�  9� }���z  �z 	�z 	B ���z 9�� :n �p�:� 	~���3  �7  �3 	�7 	B ��`   � �:� �@�(|�bX  b�  ��� �9��`�(|�ct  a�  ����;_�9�� :�%�p��:  �z � �7  �w � :���:_� ;21ِ�;  		�b�  c;  �  ��  � 	�� 	B ������b�Afzt������ �y� "� �;`�i~�ڪ-�  z��}��@� :1 ψ�:  ��  �_��zn�;  	�;|0����;  �.  �; 	�. 	B ���� �� ������r�_���_�:� p��:� � ;  �  � b�  8�p8�  D  �7  �w �� �:  �z ��    H
��}�[0�:9� 	}����  ��  �� 	�� 	B ��`   `   �} �:S�� �(|�b  bW  ���� �:� � �(|�b:  b�  �_��:��P9�@@Q�y� b�  ��  �� ;?��:y>�Ȉ�S  � � �U  `   �� �:�� �(|�c  b�  ��� �;t0�@�(|��_��9�� 9�@@Q΀y� ;  )���  �� 	�� 	B ���� �� �� :�P:_� �  �� �� ��  :��P; @@S�{ b�  :  ~	��  � 	� 	B ��� � � :� D�t  �v  ;_� ;?�P9� Fy���:`  A� 4}����  �  ~7�@@� DB@ �� 	� 	~7�@A��@� ,:` y�aN   A� ~I�~���~���:s ~7�@A��:  @� :   
  z ��c �?얊��) �@� ��} �:�H���(|�   I��6�A�[�1 
a�  b�  ����� �:N`� �(|�c6  bW  �����_���A���z:���� �{ "�z �9��i~�z�-�  {N�~��@� 9� �p�;  ��4  ����z��:@ ~I�:x����0  �3  �0 	�3 	B ��� �p � �s �������������;A p��;?� �: :� ��  �� cC  8��8�  D  �`   �� �:W � �(|�b:  b[  �_�� �;8�`�(|�bn  c  ����� Fz����  z� b�  �@�Hj� ~1�| Hz��z� {z :   �P:`U}��*{Gb  cD  c  a�  K��N   9� A� 9�  
  y� p�b� �얋?�) �@� h�] �:2`���(|�b�  b;  �_��� �:wx� �(|�b  bo  ����;�H:�@@��  R���� :���5     J2T��̈�3�>�U �8  �X H (`   �= �:���`�(|�cr  b�  �_��] �:��� �(|�b  b�  ����� Fz���  { c  ���Hk {�| Hz3�z2 zr ;@  ���: �}��*z�GcC  bD  b�  a�  K��M�  9� A� 9�  
  y� p�b� �얋?�* �@� d�� �;v�� �(|�c  cq  ���} �;S��@�(|�bV  cW  ����9��H9�@@��  Q΀�� :���  �4 ��  �/ `   �} �;� �(|�b2  c  �_�� �;P(���(|�b�  cU  ����:�� 9�%ΰ�� &{/��o  �/ �. �n  :� :_� :4А��S  �� �� �P  :��0:�� :�C֠���@�  �5 �6 �  9��@:?� ;qRۈ��O  �� �[  �� ;_�H:��    K1�6�@ZAV$2�};4]٠��  �: �  �9 ����������z����� �z� "� �: �i~ߊ�-6  zT�~�@� :� נ�;  ғ  ����z��:� ~��:\@����  �  � 	� 	B ���� �� ��������������:� p��;� � :@ �T  �T b�  8��8�  D  ��� &z���  �N �Q �  �  �� �� ��  ��@��  �� �� ��  �[  � �O  � �9  � �:  � `   � �:t	���(|�b�  bu  ����� �:�	0�`�(|�cn  b�  ����:_� ; @@S�{ ;  )��  � 	� 	B ��� � � :?� �^ Vzp�;@ I���  ��  �� 	�� 	B ���� �� �� �� :��P;`@@S{�{{ b�  9� }���o  �o 	�o 	B ��   L%��@����T��o �o �o ;< 4�  �  :_� :�P;@ F{V��:   A� 4~���  �  }��@@� DB@ � 	� 	}��@A��@� ,:  {QaM�  A� ~)�~���~���: }��@A��9� A� 9�  
  y� p�co ��얋?�* �@� �� �:�	H���(|�����] �::	`ꀁ(|�b�  b3  �_���������A�{p������ �y� "�� �; �iʪ-8  z�~��@� :� װ�:  ��7  �_��zu�:� ~��;\	x����z  �u  �z 	�u 	B ���� �� �� �� ����������:� p��:�� �� :@ �V  �V b�  8��8�  D  �`   �} �:�
(�`�(|�cn  b�  ����] �:�
@� �(|�c0  b�  ���;� :�@@R��z� :@ ~I���  �� 	�� 	   Mso����@o���B ���� �� �� :�� �^ Vzt�;` i���  ��  �� 	�� 	B ���� �T �� �V :��P; @@S9�{9 b�  :  ~	��1  �1 	�1 	B ���1 �1 �1 :�
X�  �W �w �  �U �u ;� 9��P:� Fz���;@  A� 4}����  �  }��@@� DB@ �� 	� 	}��@A��@� ,;@ z�aM�  A� )�~�Ю~Ю;Z }��@A��:  A� :   
  z7 ��b� �얊_�* �@��} �:�
`���(|�a�  b�  ��� �:
x���(|�a�  b  �_�����z6��^ _�V �� H� z��;.p�p��� ���;
��`�{' � �x(: 	|�z�cp  c  ��:���@�zv' ꀁx(6 	|�z���_�:� p��:��;?� �� �7 9� ��     N�X���t�# y�� b�  8��8�  D  ��_���A����z.��N �_��7 ;  �  � b�  8��8�  D  �`   �� �:�ꠁ(|�b�  b�  ����} �;[(� �(|�b  cS  �_��:?�l; @@b8  �8  :� 5��  ��  `   � �:�@���(|�a�  b�  �_��� �:X�`�(|�bx  b  ���\ 6�_�n`   �� �:�p� �(|�b4  b�  ����� �;o��@�(|��_����na�  �`�Hi� 9�| Hz�z { :�  ���: �~��*z�Gb�  bD  b�  b�  K�C`t  `�  z� ��}� �y�z{y }��y�zz,: 쥛?�{8���_�*�?�:��~_�*z1Gb6  bU  ꀁHjO �`�@}�| H}��| Hb�  z�� z��z�� y�,)9  zx ��| H �   OP
�հ��*^��y�z{Z!y��z�,�_�n`   � �;t����(|�a�  cq  ���] �:�����(|�b�  b�  �����na�  ���Hi� Z�| H:�  b�  bd  K�|{�| H�9���}��x��?�� h:_��:��:��;?�; �� `�@�z�' ꀁx(. 	|�z��cN  b�  �� "�`�z�' � �x(; 	|�z3�bt  b�  �� 2�@�{/' ���x(/ 	|�y��cT  c5  �� B�`�{' ���x(1 	|�z��cn  c  �� RbC  ~��b  N�!:� ; @@S9�{9 ;@ I��3  �3 	�3 	B ���3 �3 �3 ��� Vz4�-�  z��~Ԫ@� ; ���;� ��  ��  9��P:@@@RR�zR a�  ;@ I��W  �W 	�W 	B ���W �W �W ;< C�y  �n  :� :?�P   P���}�5�⎍;  F{��:�  A� 4~����  ��  ~6x@@� DB@ �� 	�� 	~6x@A��@� ,:� {aN   A� i�~Р�}�:� ~6x@A��;@ A� ;@  
  {R ЈbW ��얋?�) �@� H �`   �} �9��ꠁ(|�b�  a�  �_�� �9�� �(|�b6  a�  ���⢟�nb�  �@�Hj� 9�| H:`  bc  b  K�|n�| H�:���~�������] h;��9��:<�:��:� �] `� �y�' �`�x(4 	|�zy�c4  a�  �� "� �z.' �`�x(. 	|�{p�� 2�`�z�' � �x(/ 	|�{3�bt  b�  �� B���z�' � �x(; 	|�z.sa�  b�  �� Rc  ~I�cB  N�!:� 9�@@Q�y� ;  )���  �� 	�� 	B ���� �� �� ���   Q�?�N���>(���^ Vz{�-�  {v�~;�@� :� Ѱ�9�� ��  ��  :��P; @@S�{ b�  ;  )��  � 	� 	B ��� � � 9� 4�  �  :_� :�P:� Fz���;`  A� 4~���2  �  ~1�@@� DB@ �2 	� 	~1�@A��@� ,;` z�aN   A� }��~2خ~�خ;{ ~1�@A��;  A� ;   
  {8 Ȉc �_얉��) �@� AՀ#K���`   � �:�(���(|�b�  b�  �_��� �9�@ꠁ(|�b�  a�  ���;��; @@S9�{9 cx  ;@ I��8  �8 	�8 	B ���8 �8 �8 �8 �� Vy��:� ~��cs  �T  �S  �T 	�S 	B ���� �� �� �� :; F�؈� �z:�� �z8' ���x{0�(8 	|�yЃ�������y��z��:���   R�93&#�y��]�x:R Ԑ����z���`�z�' �@�xzv�(; 	|�{V�b�  b�  ���4  )� @A� DA� @:������y��~7��@�  z�' )2 	@� z' )� 	@� ~7�@AՀ#@��tH  D�_��z{�;[ �؈���{Y�� �{T' � �x{�(4 	|�z6�b�  cO  ���������:����z��~p�P~{�����;< C;   ~9��Ȉ�Q  �R  �� Vy��b�  :�@@Rրz� :� ~����  �� 	�� 	B ���� �� �� �^ Vz{�;  	��0  �;  �0 	�; 	B ���0 �P �; �[ `   �� �9�Xꀁ(|�b�  a�  ���� �:Up�`�(|�bx  bY  ���:��: @@R1�z1 b  ;` i��:  �: 	�: 	B ���: �: �: �: �� Vy��:� ~��b  �     S�
&��h]FN��  � 	�� 	B ���T �t �V �v ;0 Fـ�� �{;�� �{:' ���xz8�(: 	|�y���������y��z��:���:� Ԩ��@�z�����z�' �`�xzғ(0 	|�{r�bP  b�  ���T  ) @A� DA� @;?������y��}�Ȁ@�  {' *7 	@� {5' )5 	@� }��@AՀ#@��tH  D�_��zv�;v ۰�� �{p�ꀁ{z' ���xz��(: 	|�yыb.  co  ����������:����{2�~u�P~p�����:��p;@  t�۠��;  �2  9���9�@@Q΀y� a�  :� ~����  �� 	�� 	B ���� �� �� ;  	��5  �/  �5 	�/ 	B ���u � �U �o � �O `   � �;t�� �(|�b6  cw  ����] �9��� �(|�c     T���TחY0��8a�  �������{3�:   S�ژ�9�  c[  ��  �� �� �� :  �:  :�����z�' ���x(2 	|�yֳ�� ":��ꀁz�' � �x(8 	|�{4��� 2:  � :� 9��Ϙ��`�{Q��@�{N' ���xz[�(. 	|�z��cx  cY  � �� x:���:���:�p�} p� �z�' ���x(2 	|�yыb:  b�  �U "���z' � �x(9 	|�{�b�  b  �� 2b�  ~i�b�  N�!`r  :��t:   t�۠��[  `   �] �;:�� �(|���� �:�����(|�a�  b�  ����9��t:`  ~Κ�p��6 b#  K��`r  �_�z[��옃_옣?�{Y�c8  � �Hk7 ~��| H9�   �z�'y� y�zz� ���:��~<�*y�Gb�  bd  a�  b&  K��   Ux�Qmý�R]4wN   :@ @� :@  
  z[ ��cz �_얊�) �@� ��� �;7�� �(|����� �:����(|�b�  b�  �_������"�A&{t������ �y� "�� �; �iʪ-�  z��}��@� :� Ϩ�:� ���  �_��zq�:  ~	�;\(����z  �q  �z 	�q 	B ���� �� �� �� ����2������:� p��9�� �� :@ �V  �V b�  8�08�  D  �`   �} �:��`�(|�cv  b  ����] �9��� �(|�b8  a�  ���:�� :�@@R��z� 9� }����  �� 	�� 	B ���� �� �� :_� �^ f{s��  �� �� �� �3 �� �2 �  �� �� ;?�P; @@S�{ c/  :� ~���  � 	� 	B ��� � � :� 4   V
er�6����U  �Y  ;� :�P9� Fy���:   A� 4~)���  ��  ~7�@@� DB@ �� 	�� 	~7�@A��@� ,:  y�aN   A� ~I�~���~Ӏ�: ~7�@A��:� A� :�  
  z� ��c ��얊��) �@� ��] �;:�� �(|�b2  c3  �_��� �:����(|�b�  b�  �_��������B�Fz����� �{ "�0 �: �i~��-�  z�~P�@� :� Ұ�:� ���  �_��{o�9� }��:�(����  ��  � 	�� 	B ��� � ����R�����:� p��:� �v :� ��  �� b�  8�P8�  D  �`   �] �;R��`�(|�ct  cU  ����� �9��� �(|�c0  a�  ���;� :`@@Rs�zs :� ~���x  �x 	�x 	B ���x �x �x    W����Y��)�hV�:�� �^ f{r��  � �� �� �2 �� �6 ��  �� �� :?�P: @@R�z b7  :` ~i��  � 	� 	B ��� � � ; �X  �x �Q  �q :_� 9��P;  F{5��:�  A� 4~����  ��  ~.�@@� DB@ �� 	�� 	~.�@A��@� ,:� {3aN   A� ~i�}Ҡ�~Ϡ�:� ~.�@A��:  A� :   
  z ��b� �얋_�) �@� ��} �:;ꠁ(|�b�  b9  ���} �:� ���(|�a�  b�  �_���� fz��a�  :@@@RR�zR �N  �N �N �N �N � fz5�� &{3���  �s �u ��  `   �] �:�8���(|�b�  b�  ��� �:TP���(|�a�  bY  ���:�\;`@@S{�bo  �o  :���;U�ڨ���  ��     X_bV���qV��`   �� �:7h� �(|���� �:T����(|�a�  bY  ���;�`9�@@Q�cu  ��  ;_��:���Ј�v  �{  `   �� �:7�� �(|���� �:T����(|�a�  bY  ���9��l:�@@a�  ��  :���v  �o  `   �} �:��� �(|�b8  b�  ��� �:���@�(|�bN  b�  ����:���;_� :�%�Ј�u  �u �v �v  ����b�f{7���� �z� "�W �9��i}�z�-�  z��Wr@� ;{ �؈:` f�z  ���z8�;  )�:������T  �X  �T 	�X 	B ���� �t �� �x �_���Ar�����9� p��:�� �� ;@ �N  �N a�  8�p8�  D  ��6  �� �� �5  `   �� �;o`� �(|�c  cs  �_��= �:x   Y��,��\��W�Y���(|�b�  b  ���;_�9�@@Q΀y� cV  ��  �� :�8��  ��  9���;`  ~o��x�:Z �Ј�3  � � �2  :��; @@S9�{9 b�  �8  �8 ��  �� �� ��  `   � �:���`�(|�cn  b�  ����} �:�� �(|�b8  b  ���:_�;_� :�%�Ј��  �� �� ��  �������A�{o������ �y� "�o �: �i~?��.1  y��/�@� ; ���:� r��  ���z��;` i�9������n  �z  �n 	�z 	B ��� � ������������; p��:�� �� ;  �8  �8 c  8��8�  D  ��  �� �� ��  H ܋�m)  A� T�} X;_��:?�m� P���z.' ���x(. 	|�z�{a�  b9  � "��_�� B   ZlT��r^���8�  cC  ~	�bb  N�!�� �:V8�`�(|�cv  bW  ����� �:.P���(|�a�  b9  ���:��:�� ;T%ڠ��  �u �z �  ���������z2����r �{n "�� �9��i?z�-�  zT��@� :� ؠ�:` r�x  ����z��:  ~)�;|h�����  ��  �� 	�� 	B ���� �� ������_���_�:� p��:�� �� :� ��  �� b�  8��8�  D  ��:  �� �� �5  H \`   ��m*  A� T�� X:��;?�m� P�`�{2' ���x(2 	|�zӛbv  c7  �� "��_�� B8�  b  	�a�  N�!�] �9��� �(|�b:  a�  �_��] �;2��`�(|�bv  c7  �������������y����� �{ "�0 �;`�i_ڪ-:  z�   [f�-뚊x�XC�~P�@� ;9 �Ȉ:` ��r  ����z��:� ~��9������  ��  �� 	�� 	B ��� �. � �5 �_���A������: p��:� �p :@ �P  �P b  8��8�  D  �`   �� �:��ꀁ(|�b�  b�  ����= �:���`�(|�cx  b�  ���;_�l:`@@cR  �r  :���  ��  `   �� �:�����(|�a�  b�  ���� �:� �`�(|�cx  b�  ���:� :S%Ҙ��� &z���  �� �� ��  :?� :� 9�4΀��  �q �n ��  ;?�0;� :xC�����  �� �� ��  ;_�@�A@9�� :�R�x��  �z �  �t :��H;� :�]�����  �� ��  �� :�;� ;h�؈��  �� �� ��  �_���A��A�{o�����   \�(/[+�~���� �z� "�O �;`�i~�ڪ-�  y��O�@� ;{ �؈;`o�z  �_��{v�9� ,}��;\����z  �v  �z 	�v 	B ���� �z �Z �� �v �V �_���A��_���_�9� p��:�� �� ;` �o  �o a�  8��8�  D  ��^ &{v���  �R �V ��  �n  �N �Q �q  �S  �� �� �Y  ��  �� �A@��  �� �W  �w �U  �u �8  �x �p �0  `   �� �;/�ꀁ(|�b�  c7  ����� �;N��@�(|�bT  cU  ����;� ; @@S�{ cs  :  ~)��  � 	� 	B ��� � �� Vy��;  )�cw  ��  ��  �� 	�� 	B ���P �P �W �W :� F�؈ꀁz��� �z�' ���x{�(3 	|�yԣ��������y��   ]��KrW�]��z{6�:��:� а��@�z����z' � �xz��(; 	|�z:�cR  b  �_��  * @A� DA� @:�� ����y��}4��@�  z�' )� 	@� z�' *6 	@� }4�@AՀ#@��tH  D����z��:; �؈�@�z3��@�z0' � �xzZ�(0 	|�{�cN  b/  ��������:�� ��z��u�Ps�؈��� fz2�;@  }��ϐ���  �/ � �� �� �� �� ��  �4 � ��:{ ~p�����:?�;@@@SZ�{Z b2  9� }���R  �R 	�R 	B �����z�  ��b#  b�  b�  K�C-�  z9�}Ѳ@� ;9 �Ȉ� �y���`�y�' � �x{x�(3 	|�z�c  a�  ��������y��{R�:���:R א�� �z��� �z�' �`�xz9�   ^i ~a3��م��<(; 	|�zy�c4  b�  ����  * @A� DA� @;�����y��}:��@�  {R' )� 	@� {' *6 	@� }:�@AՀ#@��tH  D���z;�:{ �؈� �zu�ꀁzw' ���xz��(7 	|�y��c.  bo  ��������:_��A{v��P������:��:�  ~t�Ӡ��3  �6  9�� 9�@@Q΀y� a�  :  ~	���  �� 	�� 	B ���� �� ;@ I��r  �o  �r 	�o 	B ��� � `   � �:��ꀁ(|�b�  b�  �_��= �:��� �(|�b  b�  �_�����z.�� /�� ;�����y���`�{' � �x(2 	|�{3�bz  c  �W :��\���z5�ꀁz�' ���x(. 	|�y��b�  b�  � ":_�`�_��{s����zP' � �x(0 	   _u>5������|�z7�b�  bO  �� 2:�� ���{4�ꠁz�' �`�x(: 	|�{u�b�  b�  � B����z���� �� R�_��zx��^ ��X b���{5�� �� r����z���� ��� ��_��z{�� �� ����z:�� ��� �����z���^ ��O ����{.��^ ��N ����z5��� ��� ��_��zt����� �� H�X {y�:p�Ȉ�� ��":<�ꠁz2' �`�x(2 	|�zu�b�  b/  ���:����@�z�' �`�x(8 	|�{z�cX  b�  ��: p��:����H:�� ��@�� �� :@ �P  �P b  8� 8�  D  ��_���A2���z���� y�����{:��Z zt�����y��� &{1��_��zz��� 6y���_��zu��� Fy���_��zz��� Vy���_��zn��N f   `��2�J�b�jzz�����y���� vy������y���� �y����P����y���� �y����X����y���� �y����`����y���� �y����h����y���� �y����p����y���� �y����x����y���� �����@���xy�����y�' ���xy�(7 	|�zғbV  a�  ��������py�����y�' �@�xz�{(6 	|�zO{a�  a�  ���"�@���hy�����y�' ���xz�(6 	|�y�bV  a�  ���2�����`y�����y�' �@�xz�{(6 	|�zO{a�  a�  ���B�@���Xy�����y�' ���xz�(6 	|�y�bV  a�  ���R�����Py�����y�' �@�xz�{(6 	|�zO{a�  a�  ���b�@�zn����zw' ���xy�(7 	|�zғ�_�r���   a�1j?�U���({O����{V' �`�xz�s(6 	|�znsa�  cW  ����@�z���`�z�' ���xzr�(: 	|�yғbV  b�  ������{3��@�{.' ꠁx{O{(. 	|�z�{a�  c7  ����@�{��@�{' ꠁx{R�(. 	|�z��bN  c  ���� �z7����z3' �@�xz��(3 	|�{Y�c.  b/  ����ꠁz���@�z�' ���xzU�(7 	|�zիb�  b�  �_���@�{q�� �{o' ���x{:�(/ 	|�y���_��;��:���:���:��:��:�:_�:?�p;?�`9��P9��@;�0;_� � �� �� ��  �� (�p 0�P 8�0 @�0 H�� P�� X�p `�P h��H�� p��@�� x;  �  � b  8�08�  D  �`   � �:���`�(|�bp  b�  ���] �;2�   b�6��w�v^^��y���(|�a�  c;  �_��9��:�� :�%ָ��  �� �� �  �����B�AFzq���� �z "�1 �9��iz�-�  z7�Q�@� :� ڸ�;  p�  ���z��:` ~i�:�����0  �2  �0 	�2 	B ���_���AR�����9� p��:�� �� ;  �  � a�  8�P8�  D  ��  �� �� ��  `   �} �:SP� �(|�c:  b[  �_��= �:h���(|�b�  b  ���������b�Afzx������ �z� "�8 �;`�i_ڪ.:  {�~8�@� : р�:� P��  ����y��:� 	~��:\�����r  �u  �r 	�u 	B ������r�_���_�:� p��:� � :� ��  �� b�  8�p8�  D  �`   �= �9�����(|�a�  a�  ���   cZ'��� �);�n<�} �:S�� �(|�c:  b[  �_��;� : @@R�z c  �  � � � :� �6  �� �� �8  9� 
���ꠁy���`�y�' � �xzu�(2 	|�{5�b�  a�  �_������z��z�:0��9� �p�� �z4��`�z2' � �xzx�(2 	|�{8�c  b/  ���⊱  ) @A� DA� @;� ����z��}�؀@�  {P' *0 	@� {t' )4 	@� }��@AՀ#@��tH  D�_��zy�; �Ȉ���{�� �{' ���xz/{(5 	|�z�{a�  c  �����_���A�:� �A�zt�0�P.�Ȉ:. ~5�������� &y��:�  ~غ���;t ۠��V  �V �[ �[  ��;3 
1�Ȉ�?�:�� 9�@@Q΀y� b�  ��  �� �� �� ��  ���z�     d�Ch�:A&R0���b�  b  c  K�C.7  z��~��@� :� ԰��@�z���`�z�' � �x{r�(3 	|�{2�bP  b�  �������y��{�:���:� װ�ꠁz���`�z�' � �x{u�(3 	|�{5�b�  b�  ��⊗  ) @A� DA� @:_� ����y��}���@�  {' *6 	@� zZ' ): 	@� }��@AՀ#@��tH  D�_��{s�;3 ٘�ꠁ{1�� �{7' ꀁxz�(7 	|�z��b�  c/  �����_���A�:�� �A�zx�~6�P~0���:� ~�������;<:�  }���Ȉ9� ����o  �O �O �N �N �n  ��:3 ~0�����:��P:�@@R��z� b�  ;  )���  �� 	�� 	B ���� �� 
��{  ��b�  b�  a�  K�C.8  z��W�   e[$�K���)EQ�@� :R ڐ��`�{N��`�{Q' � �xz{�(1 	|�z�cx  cY  ������z��z��:V��9� �x����zN��`�zQ' � �xzw�(1 	|�z�b�  b[  �_��2  ) @A� DA� @;�P���z��}���@�  z�' */ 	@� {' ). 	@� }��@AՀ#@��tH  D�_��zq�: Ј����z��@�z' ꀁx{W�(9 	|�z��b�  b  �����������;�P�A�zv�~8�P~;���;[ Y�Ј�?�� Vz��:�  }�π�9� ΰ�:@ ~I��o  �n  �o 	�n 	B ���/ �o �. �n �_�;: F4�Ȉ���:���:�@@R��z� b�  :� ~����  �� 	�� 	B ���� �_�zS  ��b�  c  be  K�C.2  z��}��@� :1 ψ�   f�´mxE0?xSkJ�`�y���@�y�' ꀁx{[�(9 	|�z��cv  a�  �����_��zp�z�:0��; ���ꠁz.��@�z9' ꀁx{U�(9 	|�z��b�  b/  ����q  ) @A� DA� @:����_��zv�}���@�  z�' *0 	@� z�' )8 	@� }��@AՀ#@��tH  D���{:�:� �Јꠁz�����z�' �`�xyի(1 	|�{u�b�  b�  �_���������:����{:�}��P}��x����� fz��;`  ~q�ӈ��S  �� �� � �3 � �: �Z  �� �� ���9� }��p����:��P;`@@S{�{{ b�  :` ~i��q  �q 	�q 	B ���q �q ��{  ��b�  b  c%  K�C.8  z��~U�@� :� Ҹ����zZ����zN' ꀁxy��(. 	|�   gm��b� w'Zoz��b�  b[  �_���_��zq�z0�;1��: ـ����{8�ꠁ{/' ���xz��(/ 	|�y׻b�  c;  �_�⊙  ) @A� DA� @:��P�_��zq�}���@�  z0' *0 	@� z�' )8 	@� }��@AՀ#@��tH  D���z��9� �x����y���@�y�' �@�x{W�(9 	|�zW�b�  a�  �_�������;�P��z��}��P}��x���;\�;   }���Ј��  ��  :� :S%Ҙ�:  ~)��  �  � 	� 	B ���� �� �� �� ��������A�{y������ �z� "�� �:`�i~?��.1  {8�~�@� ; ���:� ���  ���z��9� }��9� ����N  �R  �N 	�R 	B ���_���A��������:a p��;� � :  �3  �3 bc  8��   h��L��ui��N_�8�  D  �<Ȃ̂�Ђ�ԁ�آ\ܑ��
�_��?�����������H �`   �� �;n��@�(|��_��� �:��� �(|�c  b�  ����) �@� ��� �:O� �(|�c4  bU  ����� �;n(�@�(|��_�����������z8����x �zo "�� �:@�i?��-�  {�~��@� :� ՠ�9� z��  �_��{w�:� ~��:@����0  �7  �0 	�7 	B ���p �w �����������:A p��:�� �� :� ��  �� bC  8� 8�  D  �`   �] �;z����(|�b�  cq  ���} �:�����(|�a�  b�  ���9� ���`   � �:���@�(|�bZ  b�  �_��� �:6� �(|�����} H�� z��;/p�x�� ��; ���   i�6)D��>(�T�{' �`�x(2 	|�{nsa�  c  ��;_�����{S' ���x(3 	|�z��b�  cO  ���;! p��:��:�� �� �� :@ �Y  �Y c#  8�8�  D  ��_���A"���z8��X zw�����y���V {p��_��zq��� &y���_��{v��V 6zn��_��{q��Q Fzo��_��{v��V Vzq��_��{r��R o�_����z3��@�z;' �@�xzV�(; 	|�{V�b�  b3  �_��`�y��� �y�' �`�xz;�(6 	|�z{�cr  a�  �_�"�@�y�����y�' �`�xz��(/ 	|�{z�cR  a�  �_�2� �{����{' ���xy�(; 	|�yыb2  c  �_�B�@�z����z' ���xy��(; 	|�y��cR  b  �_�R� �z�����z�' �`�xz��(/ 	   jgd�r5��ѮEr|�{x�c  b�  �_�b9��`:�P;_�@:?�0:�� �� � �Y �9  �� (�� 0�� 89� ��  �� c#  8� 8�  D  �|�������|Ă\ȡ�̒_�
��������������H  TAՀ#��| Hb:  ���� �  ��~��N� AՀ#����| Ha�  �\��y ��  ؈~��N� � H�X zq�:�Ј�� ��2�������;A p��:�� �� ;  �:  �: cC  8�08�  D  �A݁�8!�� (|�����N� !        ������� u�      ���         T   H �       H    ��� �                   ,        0@  7    07         ��� `       T   H �       [�       k7��zP�͐�،��� ��                   0      �  4   �7    �7    �7    <7    p7    �  � H     h7    x  t L     T     �7    �7    �7    	@7    	`6    	�7    
�7    47    �     �7    l7    �7    �7    �     �7    $7    $7    �     �     7    �7    �7    7    ,6    `7     7    p     x     7    $6    `7    �     ,     4          T     \     7    @7    `7    �7    �7    �7    6    H7    0     8       l�݈jZ~��� �7    �6     7    !�     !�     ",7    "�7    #�     $#     $l     $t     $�#     $�#     %     %     %      %,     &D7    '     '     '�     '�     '�     '�     (�7    )�     )�     *d7    *�7    +07    +�     +�7    ,�7    -7    -�7    -�     -�7    .�7    /,7    /�7    0$7    0`     0�     0�     1<7    1\6    1�7    3      3(     3�7    3�6    47    5�     5�     6�7    6�7    7�7    7�7    86    8@7    8�7    8�7    9x7    9�7      m1d�r��1/q 9�6    :7    :�7    ;H7    ;h6    ;�7    <�7    <�6    =7    =�7    =�7    >7    >87    >X7    >x7    >�7    >�6    ?,7    @l7    @�7    A87    A�     A�7    A�     B     B<7    B�7    C7    C`     Ct7    E�7    E�7    J�7    K7    K06    K\7    L7    L,6    LX7    L�7    M@7    M�7    N     N(     N@7    NH7    Nh     N�     N�7    O7    O�7    O�     O�     P7    P7    P<     P�     P�7    P�7    Q|7    Q�     Q�     Q�7    Q�7      n��Ǽ%Tz""� R4     Rt     R�7    R�7    Sp7    S�     S�7    T     TT     T|7    T�7    UP7    U�     U�7    U�7    V47    VT6    V�7    W�7    W�6    W�7    X�7    X�7    [<  [8 [P"    [d  [` [x"    [�7    [�7        ��� ��       T   H �       h    ��� �0                   ,        0 `   �7    7    P7         ��� �`       T   H �         �    ��� ��                   (        ,     H7     p7             D D        8       D � 	d 
   oȞAȊ��#���� 9l :T [P [T [x [| [�    h             	                	                            	                        @                         �                                U                              �                             �                        ���          �                        :X     �                  1A    ���          �                        ;�     �                        ���          �    �               p�i�i�C�v]�           �                                      �                                                                                }                      ����                                        � �                              �                                   @ �� �                           �                                   @ �� K                                                       ��������        �A���a�����|�� (�!�A`]  �A  < D� �a `3� `   qm��Ċ�����X| �A݀`~  � `� `��m)  A� \� X;���A `�Z `;:m� P���{6' ꠁx(6 	|�z��b�  c5  �� "��_�� B8�  cc  	�c�  N�!;>  ���� /�� ��A `�� `�A ��W�� ���:�
@;�  b�  :� ~����  �� 	�� 	B ���^ /�V ;  �6 0;  �� A�� H� z��;|����� � ��@�z�' ���x(4 	|�z��cT  b�  ����;� p��;���| ;  �<  �< c�  8� �8�  D  � @)� �@� \�� �;_��� `� `;t��= �뀁{v' � �x(6 	|�{�c�  cu  �� ":�  �� 0�� 8cC  )�b�  N�!� `�x `;�
@�� @* �@� \� �:����A `�: `:��� ��`�z�' ꠁx(< 	|�z��cr  b�  �V "   r�>FA�A>�D"C;@  �V 0�V 8b�  	�b�  N�!A݁�8!�� (|��A��N� !        ������� |�          < d 	    �� �!�(�A�3|�� (�!��`]  �A  < D� 3�  | �A݀`~  � H�\ {z�;���Ј�\ �A r�^ &{|��\ &{z�� ���;� `��;���| ;@ �\  �\ c�  8� p8�  D  �A݁�8!`� (|���#N� !    ������� }`          8  � 	               @           ��� �    ��                                         be< 
�be< �be< V be< Y�be< Z be< i�        be< � be<  �                        �  ��                     s
I�j�f�u       ���  ��� �        ��� ��0�}�� 4p0�}�� 5�        ��� ��0�}�� 3���� �@��� ��        ��� � 0�}��  ��� ~���� ~                                 �              �    �    ��� �         R�haG��                        �#�G��aF        ��� ����� �P                                                                                                                                                                                                                                           t���%ڢ���  P                  X    ���  ��� � ���  ��� }�                                                          `                            C��       \     ��� `��� � ��� `��� }�0�}�� 0 0�}�� 2�be<                                     �                            ��{� �     x    ��� ����� � ��� ����� �H                                                          �   n   +                      K�E  �      �    ��� �`��� � ��� �`��� �                    u5�*['y�9�                                          `   6                         t�z�  �                          p��� u`                                                                  @                 ��� u�                                                                                      x��� |�                                                                   `                   p��� }`                                                                                                          v�E����t�aW�         3                                                                          ��� 0��� ���� ���� �                                        ��� � �ڜ�&��     ��                             0                                                                                                                                �   �   be< ��        be< ��        be< ؐ                         00`@00 
 %��������@@@@@@@@@@@@@@@@@@@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@                  w�[�:�߾2���    0                                           �  (          �   z               h     [\       �     [4       �     �       �     �       �     �       �     	�       �     l           	�      �     	�      �     
`      �     
d           
�            
�      8     H      P     P      h     �      �     �      �     �      �     �      �     $            (           �      0     �      H     �      p     �      �     @      �     D   xY9�`�io���O0      �     �      �     �      �     8            <           �      �     �            4           8      0     �      H     �      `     �            �      8     �      `     L      x     �      �     �      �     �      �     t      �     �           �      (     �      	     �      	0      @      	H     P      	`      @      
(      D      
@     "�      
`     !�      
x     "�           "�      (     #D      @     #H   yBO4��Ź^�l      X     #�      p     #�      �     $�      �     $�      �     '4      �     '8           )�      (     )�      @     ,      X     ,      p     .l      �     .p      �     /�      �     /�      �     1�      �     0�           1�      �     1�      �     40      �     3@           40      �     44      �     6<           5�            6<      8     6@      P     6�      h     6�      �     6�      �     7       �     7L      �     7P   z�a��
̩�O      �     8x      `     8|      x     90      �     94      �     :T      8     :�      P     ;�      �     <8      �     =0      �     =4      �     =�      �     =�            ?�      �     ?�      �     C�      �     C�      �     Jx      �     J|      �     K�      P     K�      h     L�      �     L�      �     V�      �     V�      �     X           W      (     X      �     X      �     XH      �     XL           [   �   {           {Q�[Wl��U��       p              �              �              �              �              �                                        �             �             �                          (             @             X             p             �             �             �             �                                        8             P             x             �             �             �             �             �                                     |��M�򸏧��       �                                        8             P             h             (             @             h             �             �             �             �             �                          0             	              	8             	P             	h             
0             
H             
h             
�                          0             H             `             x             �             �             �          }�xT����3��B�                                 0             H             `             x             �             �             �             �                                        �             �                                        �             �                          (             @             X             p             �             �             �             �             �             h             �             �             �          ~��;��Vc�m�H      @             X             �                           �             �             �                          �             �             �             �             �             �             X             p             �             �             �                                        0             �             �             �                          �                           �                                                          ��˾|)/:#߈                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo      "  �  ���        0�}��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ��r�'+��&9 �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ��s�Xo   `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ��s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ��s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ��s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ��s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ��s�Xo                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��s�Xo       �                                            �\@��@@@@@@@@@@a\���              �          d    ��� t���� `  E�    ��� t���� `  E�    ���   ��� `  �    ���  T��� `  �    ���  X��� `  �    ��� #X��� `  �    ��� !���� `  �    ��� #T��� `  �      �    ��������    ��    �        
     P������ņ    ���ـ    �        
     P���ن    ��ـ    �       #      P�����ً       F��� #\��� `      ��� #���� `  |    ��� #���� `   ��Q����S<�*  |    ��� $8��� `  �    ��� $<��� `  �    ��� $���� `  D    ��� $���� `  �    ��� &��� `             ��  ��� &��� `      ��� '<��� `  p      
     K������ '@��� `  p    ��� '���� `  �    ��� '���� `  �    ��� '���� `  8    ��� '���� `  8    ��� ,0��� `  d      y��������@@\����@@@@@ 	��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ �\����@@@@@@@@@@@@@@@@@��������@@@   ��@��]:�]�t/@@@@@@@@@@@@@@@@@@@@@  80����@@@@@@�������   ���� 	�  �  F���  g������  
�  �  d \����     ��� ,4��� `  d    ��� ,���� `  �    ��� ,���� `  �    ��� 0 ��� `  �    ��� .��� `  ,    ��� .���� `  �    ��� .���� `  �    ��� 0��� `  X      ��    	��������ǆ    ����Ā    �             P����Ć    ���ƀ    �    ������ǆ    �������    �        P     P�������    ������ŀ    �    \�����ŋ           ��� 0$��� `  �       ������*T4T����� 0���� `  L    ��� 0���� `  L    ��� 2���� `  �    ��� 1���� `  L    ��� 2���� `  �      L�    	��������ǆ    ����Ā    �    ��������    ���ƀ    �    ������ǆ    �������    �    ◖��@��@���@\���    ������ŀ    �    \�����ŋ        ��� 2���� `  �    ��� 4��� `   l                  ��� 3���� `  �    ��� 4��� `  �    \����   ��� 4��� `   l    ��� 54��� `  !4                   ��� 4���� `   l    ��� 54��� `   ��) �4�3gp  !4    \����   ��� 58��� `  !4    ��� 7,��� `  #�      !4�    ���������    ���ŀ    �        
     P���ņ    ��   T �    L �        
     P������Œ       # 
     P���ْ       2      P�����ن    �����ـ    �       =      P������ً           ��� 70��� `  #�    ��� 9���� `  %�    ��� 8���� `  #�    ��� 9���� `  %�      #��    	��������ǆ    ����Ā    �    ��������    ���ƀ    �    ������ǆ    �������   ! �    ׁ�������@�������@��������     �ף���BE���8  ������ŀ    �    \�����ŋ        ��� 9���� `  %�    ��� <L��� `  &�    \������ ��� ;4��� `  %�    ��� <L��� `  &�      ��������@@\����@@@@@  d\����@@@@@@@@@@@@@@@@@��������@@@@@@@@@@@@@@@@@@@@@@@@  %� 0����@@@@@@@@@����@@@���� �  F \������� <P��� `  &�    ��� <���� `  '    ��� <���� `  '    ��� <���� `  't    ��� <���� `  '�    ��� >��� `  (<                  ��� >��� `  (<    ��� @���� `  )    P�������@@@@@@@@@@@@@@  ��� @�   ��g�<��M��s���� `  )    ��� C��� `  )�    ��� C��� `  )�    ��� Ep��� `  *0    ��� Et��� `  *�    ��� G���� `  *�    ��� G���� `  *�    ��� ID��� `  +�         e     ���� IH��� `  +�    ��� K ��� `  .|    ��� J0��� `  +�    ��� K ��� `  .|      +��    	��������ǆ    ����Ā    �    ��������    ���ƀ    �    ������ǆ    �������    �    
晖��@ׁ���    ������ŀ    �    \�����ŋ       ��� K$��� `  .|    ��� M���� `  0    ��� L�   ��s�v���N�S��� `  .|    ��� M���� `  0      .|�    	��������ǆ    ����Ā    �    ��������    ���ƀ    �    ������ǆ    �������    �    ���@����@��������    ������ŀ    �    \�����ŋ         ��� M���� `  0    ��� O���� `  2d    \����   ��� O��� `  0    ��� O���� `  2d    ��� O���� `  2d    ��� P ��� `  2�    ��� P��� `  2�    ��� P\��� `  3�    ��� P`��� `  3�    ��� P���� `  3�    ��� P���� `  3�    ��� Q���� `  4X      3�      �+��=� s�y� 	��������ӆ    �����Ӏ    �    ����ņ    �����ـ    �        	     P�������       ��� Q���� `  4X    ��� R���� `  4�    ��� R���� `  4�    ��� S���� `  5       4��    �����Ԇ    ���ŀ   " �     �    �������Ӗ    ���ӆ    ��ـ    �        
     P�����ً           ��� T��� `  5     ��� U4��� `  5       5 �    �����Ԇ    ���ŀ   " �     �    �������Ӗ    ���ӆ    ��ـ    �        
     P�����ً           ��� U���� `  5�    ��� V�   �y˰���KaN��� `  7x      5�    	��������ǆ    ����Ā    �    ��������    ���ƀ    �    ������ǆ    �������    �    ���@����@���@������    ������ŀ    �    \�����ŋ       ��� V���� `  7x    ��� V���� `  7�    ��� V���� `  7�    ��� Y ��� `  :�      7܂    ������Ɔ    ���ŀ    �        
     P���ņ    �����ŀ   " �     �    �������Ӗ    ���ӆ    ��   T �    L �        
     P������Œ       # 
     P���ْ       2      P�����ن    �����ـ    �     ��^r8淙eWQK     =      P������ن    ����ـ    �       H 
     P�����ن    ������    �    \��Ć    ������ـ    �    \���Ë      ��� Y$��� `  :�    ��� ]8��� `  ;`    ��� ]<��� `  ;`    ��� c���� `  >�      ��������@@\����@@@@@  �\����@@@@@@@@@@@@@@@@@��������@@@@@@@@@@@@@@@@@@@@@@@@  ;`#0����@@@@@@�������������� �  
�  
�  �  �  d�  �  �  �  �  �  �  �  �  �  
 \����  ��� c���� `  >�    ��� d���� `  ?H      >�    ���Ԇ    ���ŀ   "    ����i;�w?̃     �    �������Ӗ    ���ӆ    ��ـ    �        
     P�����ً     ��� d���� `  ?H    ��� e���� `  @      ?H�    �����ǆ    ���؀    �    \���؆    ����ـ    �    \��Ӌ     ��� e���� `  @    ��� p��� `  A�    ◖��@����      ���������@����    @�    	��������ǆ    ����Ā    �    ��������    ���ƀ    �    ������ǆ    �������    �   �    �     
o���������    ������ŀ    �    \���׋       A�@@@@@@@@@@         ��� p@��� `  C�    ��� qd   �JS��W`&5�.���� `  D�    ��� p|��� `  C�    ��� qd��� `  D�      C��    	��������ǆ    ����Ā    �    ��������    ���ƀ    �    ������ǆ    ������ŀ    �    \�����ŋ           ��� qh��� `  D�    ��� q���� `  E�    ��� q���� `  E�    ��� t`��� `  E�     
��������@@\����@@@@@ @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@       @@@@@@@@@@@@@@@@@@@@@@@@   \����@@@@@\����@@@@@   	\������@@@@@@@@@@@@@�   0@@@@@@@@@@@@@@@@@@@@@@@@@@@@��������@@@@@@@@@@@@@@@@@@@@@@@@@\@@@@@@@@@@@@@@@@@@@   ����cȅ����u@@@@@@@@@@@@@    @@@@@@@@@@@@@@@@@@@@@@@@@@@@ �\����@@@@@@@@@@@@@@@@@��������@@@@@@@@@@@@@@@@@@@@@@@@  E�40����@@@@@@�������������� F��g���������������� \����      ����@@@@@@@@@@         ��� `                                                                                                                                                                                                                                                                                                           �����}	K���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo       �     �  �                                               �                               �     0          @          @                                      �          @              �                                                                       �                      @                                                                                               @              �                                    �                                                      ��s�B�pI1��E              �                                                                                                  �                                                                                          @                           @         /   �          8   c    �%��}�E�q�e�-���A 	 �#)%&I&�'u'�(�)i*1*�+]./�22e3-3�3�4Y4�5�77y:5:�>�>�?�A=C1D]E%G}   �               m��m���   ��������       �������   ؃�m��������m�����   	؃�m�����   	؃�mӒ���   ����   $���mƤ������m�   ����
�~��ƈ���mŧ�������mȁ�����       �@��@��ą�����ň   �@��@���È   �@��@������������ɕ��   �@��@���ŗ����             0�}�� 4�0�}�� 5p                        0�}�� 5�                0�}�� 5�                              �   �              7   +   �      w   L   	�      {   Y   �      �   f   �     ~   �         �   �         �   �   �     �   �   �                                                                                              0�}�� 6X                                   ��>����}���                0�}�� 6�                        �ةF1�                                  h                                                                                                                                                                                                                                                                                                                                                                                                                                 ��r�py�^2�E                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ��s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ��s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ��s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ��s�Xo       p�  ���                   �      �           <   c    �%�Q�}�E�q�e�-���A 	 �#)%&I&�''u'�(�)i)�*1*�+]./�22e3-3�3�4Y4�5�77y:5:�>�>�?�A=B�C1D]E%G}                         5         	�           �     �        �                                        0             @           	  P           
  `             a             c             o             p             �             �        ���crg*�m.�'1                         �             �             
�             e             �     @         �           !  �           "  �           &  �           (  i           ,         F      -   P     F      .  �           1        �      2  �           3  
�    	      4  
�           5  
�           8              9  �            :  �           ;  �           <  �            =  �           >  �   �|)V�qs�Vs           E            +   i             j             k             r               s              t             v               x  
�           z  m           �  
�           �               �              �        �      �               �   0           �   @           �   P           �   `           �   p           �   �           �   �           �   �           �   �           �   �           �����#�7��   �   �           �   �           �   �           �              �        
      �  0     
      �  @           �  H           �  P     
      �  \           �  `           �  d           �  h           �  �           �        d      �  l           �  n           �  �     e      �  	      d      �  p           �  	p     �      �  t           �  �     	      �  �     
      �  �           �  	�     ��>�lT?��ޭ�@   P      �  �           �   �           �  �           �   �           �   �           �   �           �   �     G      �  �           �       
      �        d      �  �           �  �     h      �              �        $      �  P     k      �  �     �      �  P     �      �  
@     H     �              �             �            �             �  0          �  @          �  P          �   �\U���p�)'V�  `          �  p          �  �          $  �          %  �          &  �          '  �          (  �          )  �          B            +  G                           ��������@@@@@@@@@@@@@@@@@@@@@@�        �                                                               �                                                   M ��                           %00         
                                                                          ��v�ΜĴ��� 
                                                                                                                                                                                                                                I     H����                                               Y                     �  @                         �        � � �  	                       �   	                       �           0              �           @              �           P   �����cO��?T              �   	        `             �           p              �           q              �           s      	        �                 
        �           �              �   	        �              �           �              �                            	                   ` � �                            �                           	 @                                                                                   ` � �              �a##������           ` � �                             @	     3                  �                       `   �           u              �                                      �               �              @        � � �  	                   ` � �                          �                        �   	         p               �                        `   �                                   	                   ` � �                           	 @        y   ��%��q���=�              �                             @ �       +                             L                         F        p �                F        p �                        ` � �                           	 @                     p   �              �        p � �                      ` � �             	        � � �  	     3                 �        3   0              �   	                     `   �                             @           ��%kY�3�h           p � �                      � � �       9                  �        9                  �                       � � �       <                  �        <                  �                                                                                                                                                                                                   	    +               � � �                        `   �                                                  ��r�7�
�}���x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                          `   �                        `   �               ��{��H# -�.               	 @                   p � �        i                  �        i   
               �                            @                                                     `   �   	                     `   �   	                     `   �   	                     `   �                       � � �  	     r                   �   	     r                  �    U          r                	                   ` � �                                   3       ��?p%n��O��9              �                                     }          R   �                                                                                                                                                                                                                                                                   3   ;      #        �                      ` � �                      ` � �              �        � � �  	                     `   �   	           ��W��g�p����           ` � �   	                   ` � �   	                   ` � �   	                   ` � �   	                   ` � �   	                   ` � �   	                   ` � �   	                   ` � �   	                   ` � �   	                   ` � �   	                   ` � �   	                   ` � �   	                   ` � �   	                   ` � �   	                   ` � �                
        `   �               ��	�mډϬ�}           `   �                       `   �                F        `   �                       `   �                       `   �                       `   �                       `   �                        `   �                        `   �                        `   �                        `   �                        `   �                        `   �                
        `   �             
        p � �             
        p � �             ��3���W�%mL           p � �                     p � �             
        p � �                     p � �                     p � �                     p � �                     p � �                     p � �             d        p � �                     p � �                     p � �              e        p � �             d        p � �                     p � �             �        p � �                     p � �             ���N����#*�   	        p � �             
        p � �                                                     p � �             P        p � �                     p � �   �      �         �    t  s       �    �                      �                                       p �                  �        p   �                      p � �              
        p �                  �        p   �                �        p   �                �        p   �                ��KP���(�   �        p   �          �                                       p �                        p �            �                               G        p �     	                   ` �                              P                     `   �   	                     `   �                �        p   �                �        p   �                f        p   �              
        p �                  r        p   �    �      �         �    p  o       �   �J:�5,���    �                            r        p   �    �      �         �    r  q       �    �                            �        p   �               o        p   �              d        p �                        p �                h        p �                  p        p   �                P        p   �                      p �                $        p �                k        p �                �        p �                �        p �                  ���2#���Y�5   �        p   �                z        p   �              H        � � �  	                     `   �                        `   �                        `   �                        `   �                                                                                                                                                                                       �                                                         �                               ��&���>5��60   @                                                     �                            �                               F                         @                              7                                                        C                         �                            �                                                                                      y                                                                                     �Ybl��?NV�<�                                                                                                                                                                                                                                                                                                                                                                                                                        U                            �                     �       V                            ��S�,�-���n�   �                            �                                                                                                           #                            �                     �      $                           �                            �                     �      �                                                      �                           �                           �                            �                     �       � �գ��lZ��8  �                           u                            �                     �      v                           #                     �      *                           �                           �                           �                                                        F                           �                           �                                                        F                           �                            ���¤���gZ��@  �                           �                           �                           �                                                       �                     �                                 �                            �                     �      �                           V                           [                            f                     f      \                           �                            r                     r       ��c)��;3B���l  �                            r                     r      5                            �                     �      �                           	M                           o                    o      	N                           
�                     �      
�                            p                     p      �                            P                     P      �                     
      G                           Q                            ��Mk�D�r�q8  _                            �                     �      c                                                       z                     z      !                    �      �                           -                         �                              G                                                                                                                    '                                                            >                               ��6#���ب��                               T                           _                           ;                           8                           M                                                                                                                                            .                                                        E                 �                 �    v  w           ���`                       ���`             �           �3[�&��s��,܎         �    y  z           ���`                       ���`             }            ����      |  }           ���`                       ���`                                        �      ~         �    �               ���`                        �� #�                        �� #�                                         �      ~  �     �    �                         �                                K      �  �                            �-��,�,
_��o�                                                                                                                                           d                                                      
                                                      P                                                      	   	                           
                        �                           e                                                      ��K��硽���                  	                        �   	                   x �     	                        �              �                          �                          �                          �                      	    �                      
    �                                                     �                          �                          �                          �                          �                         ��S�E��9��    �                          �                          �                                                     �                          �               	                        �              w               	                   x �     	                   x �                �                          �               	                        �              v                          �                          �                         �H�~4�3���+FK    �                          �                                                     �                          �               	                        �   	                   x �     	                   x �     	                   x �     	                   x �     	                   x �     	                   x �                �                           �                      !    �                      "    �                      $   Ë\�8�?�,��/A    �                      %    �                                                 &    �                      '    �                      (    �                      )    �                          >                      *    �                      +    �                      -    �                      .    �                      /    �                      0    �                      2    �                      3    �                           ĉ8��1�F                         5    �                      6    �                      8    �                      9    �                      :    �                      ;    �                      <    �                      =    �                           F                      ?    �                      @    �                      A    �                      B    �                      D    �                      E    �               	             ŉ6���5������              �          F    �                      G    �                      H    �                      I    �                      J    �                      K    �                      L    �                      M    �                      O    �                      P    �                      R    �                      S    �                           G                      W    �                      X    �                      \   Ɖ�i���;J�D    �                      ]    �                                                  ^    �                      _    �                      a    �                      b    �                      c    �                      d    �                                                 f    �                      g    �                      h    �                      i    �                      k    �                      l    �                      m   ��->]�~xJ�`h    �                      n    �                          �                      o    �                      p    �                          �                      q    �                      r    �                      s    �                      t    �                      u    �                      v    �                      w    �                      x    �                      {    �                      |    �                      ~   ȩ=��J�,��28    �                          �                      �    �                      �    �                      �    �                      �    �                      �    �                      �    �                           h                      �    �                      �    �               	                        �   	                   x �     	                   x �     	                   x �     	                   x �     	           �9��Wѭ򜺊           x �     	                   x �            �    �                      �    �                      �    �                      �    �                      �    �                      �    �                                                      $                                                       k   !                        �   "                        �   #                   �    �                      �    �                      �   �О�e��:d@    �                      �    �                      �    �                      �    �                      �    �                      �    �               	                        �   	                        �               H   $            	                        �   	    +               x �                     �                            �            	                        �              9   '            	                   x �                    ��������`�  �      1   #                    4   3            5   3             �   3               3            x   3                              #                                                                !               "                                                                                                                                 	               
                        	                  ��}��Р�G��2                     (               z         
                                                                                                                                                            	      	                                          
      
                                                                        	   
                      (                        	                 ͹?��i])1  �   ����    �������      1A ����������         ����������         ���\  �    ��������    ��    �        
     P������ņ    ���ـ    �        
     P���ن    ��ـ    �       #      P�����ً              
            H       d      y��������@@\����@@@@@ 	��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ �\����@@@@@@@@@@@@@@@@@��������@@@@@@@@@@@@@@@@@@@@@@@@  80����@@@@@@�������   ���� 	�  �  F���    �0�UXB����� g������  
�  �  d \����@  ��    	��������ǆ    ����Ā    �             P����Ć    ���ƀ    �    ������ǆ    �������    �        P     P�������    ������ŀ    �    \�����ŋ     \���  L�    	��������ǆ    ����Ā    �    ��������    ���ƀ    �    ������ǆ    �������    �    ◖��@��@���@\���    ������ŀ    �    \�����ŋ                \����            \����  !4�    ���������    ���ŀ    �        
     P���ņ    ��   T �    L �          �&_%�� �2�2� 
     P������Œ       # 
     P���ْ       2      P�����ن    �����ـ    �       =      P������ً     @  #��    	��������ǆ    ����Ā    �    ��������    ���ƀ    �    ������ǆ    �������   ! �    ׁ�������@�������@��������    ������ŀ    �    \�����ŋ     \������  ��������@@\����@@@@@  d\����@@@@@@@@@@@@@@@@@��������@@@@@@@@@@@@@@@@@@@@@@@@  %� 0����@@@@@@@@@����@@@���� �  F \�����       q               P�������@@@@@@@@@@@@@@ aP�������@@@@@@@@@@@@@@ @a     e   �ִ)��9� T     �              +��    	��������ǆ    ����Ā    �    ��������    ���ƀ    �    ������ǆ    �������    �    
晖��@ׁ���    ������ŀ    �    \�����ŋ     @  .|�    	��������ǆ    ����Ā    �    ��������    ���ƀ    �    ������ǆ    �������    �    ���@����@��������    ������ŀ    �    \�����ŋ     \�����  3�    	��������ӆ    �����Ӏ    �    ����ņ    �����ـ    �        	     P�������     �  4��    �����Ԇ    ���ŀ   " �     �    �������Ӗ       у�Ф�J�O.�`����ӆ    ��ـ    �        
     P�����ً       5 �    �����Ԇ    ���ŀ   " �     �    �������Ӗ    ���ӆ    ��ـ    �        
     P�����ً       5�    	��������ǆ    ����Ā    �    ��������    ���ƀ    �    ������ǆ    �������    �    ���@����@���@������    ������ŀ    �    \�����ŋ     �  7܂    ������Ɔ    ���ŀ    �        
     P���ņ    �����ŀ   " �     �    �������Ӗ    ���ӆ    ��   T �    L �        
     P������Œ       # 
        �kOR]�$eH��uP���ْ       2      P�����ن    �����ـ    �       =      P������ن    ����ـ    �       H 
     P�����ن    ������    �    \��Ć    ������ـ    �    \���Ë     K���  ��������@@\����@@@@@  �\����@@@@@@@@@@@@@@@@@��������@@@@@@@@@@@@@@@@@@@@@@@@  ;`#0����@@@@@@�������������� �  
�  
�  �  �  d�  �  �  �  �  �  �  �  �  �  
 \����  >�    ���Ԇ    ���ŀ   " �     �    �������Ӗ    ���ӆ    ��ـ    �        
     P�����ً       ?H�       �.�
=�I�IX�%�����ǆ    ���؀    �    \���؆    ����ـ    �    \��Ӌ     ◖��@�������������@����K���  @�    	��������ǆ    ����Ā    �    ��������    ���ƀ    �    ������ǆ    �������    �   �    �     
o���������    ������ŀ    �    \���׋       A�@@@@@@@@@@         C��    	��������ǆ    ����Ā    �    ��������    ���ƀ    �    ������ǆ    ������ŀ    �    \�����ŋ      
��������@@\����@@@@@ @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@       @@@@@@@@@@@@@@@@@@@@@@@@   \����@@   ԤxVԘ]�a-c&@@@\����@@@@@   	\������@@@@@@@@@@@@@�   0@@@@@@@@@@@@@@@@@@@@@@@@@@@@��������@@@@@@@@@@@@@@@@@@@@@@@@@\@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@    @@@@@@@@@@@@@@@@@@@@@@@@@@@@ �\����@@@@@@@@@@@@@@@@@��������@@@@@@@@@@@@@@@@@@@@@@@@  E�40����@@@@@@�������������� F��g���������������� \��������@@@@@@@@@@                       �@@@@@@@@@@              �         �������    ���    ��<    �� @ ��                                                                   k             f      j  u   ռ�������[   j  {   j  �   j  �     �   #  �   a          �             c  �                           �   #   �   a   l              #   �               �     �   /      #   �        	            �      �   	            �   a   h                �       !   �      �     �   4   A         (   �                     �   !   �      �     �   4   A         (   �                  !   �      �       !   �      �      !   �      �       !   �      �   0   !   �      �Jx��.-Â��A   �   @   !   �      �   P   !   �      �   `   !   �      �   p   !   �      �   �   !   �      �   �   !   �      �   �   !   �      �   �   !   �      �   �   !   �      �   �   !   �      �   �   c                                  �   a           �       !  �   c  �                 e      f      j  u   j  {   j     g   �   g   �   g   �   g   �   g   �   g   �   g   �   g   �   g   �   g   �   g   �   g   �   g   �   g   �   g   �   o         o         !   �      �      ׯ���G�D(  �   a          
          !   �      �     �   a          
          !   �      �     �   a          
            `   #   �   !   �      �     �   a          
            a   =   ����       #   �   !   �      �     �   a          
          !   �      �     �   a          
          !   �      �     �   a          
          !   �      �     �   a          
          !   �      �     �   a          
            b   #   �   !   �      �     �   a          �N� %���..gF   
          !   �      �     �   a          
          !   �      �     �   a          
          !   �      �     �   a          
          !   �      �     �   a          
          !   �      �     �   a          
          !   �      �     �   a          
          !   �      �     �   a          
          !   �      �     �   a          
          !   �      �     �   a          
          !   �      �     �   a          
          !      #   4      ����	<*���   �   #   x     i   #   5   "   3   ;      �   L      N        �   a          
             �   #        j   #   !   !   "      �   L      N        �   a          
          !   3   %      0         �   #      !      #         �   #         �   #   
      �   #         �   #         �   #         �   #         �   #      "      }      �   L      N        �   a          
          "      �      �   L      N        �   a          
          !      #   &   �,��n��9I�   n   d   a           �         �   !           k   A                     #  �   !  �            b            �   #   s   !      #   t   j   u         a   '      �       #                    #      a           �         �         A            #   2         a   '      �       #             !   1   (   #         n  �      �         z     	            !   z     	      	   c   {                          �            j   *   l����       !  �   #   ;   ����s����mx   !  �   #   >   j   �   l����       n  �            !  �   #      !  �   #   .   !   �      �     �   a          
          !   �   !        �     �   /   L      a         	                n  �      	      !  �   #      !  �   #   .   !   ,      �      �   a   /      
          �      �     �   /   L      a         	       !   -      �      �   a   /      
       !        �     �   /   L      a         	          ,      -      M      L         �   I   �{����C���:TS   #   �      �      �                     !  �   #      !  �   #   .   "   1      !   �      �     �   /   a         	       "   1      !   �      �     �   /   a         	       "   1   #   !   �      �     �   /   a         	                       (         (   >        (   $              (   �             2            #  �   !  �            b         !   �   "   1         �     �   /   a         	       !   �   "   1         �     �   /   a   �M��XVK�*p         	       !   �   "   1   #      �     �   /   a         	                                  
      n  �   n              !  �   #      !  �   #   .   !   �      �     �   a          
          !   �      �      �     �   /   L      a         	                n  |            !  �   #      !  �   #   .   !   �      �     �   a          
          !   �      �     �   >      �     �   /   L      a         	                n  �            ��܃��%Y-��_   !  �   #      !  �   #   .   !   �      �     �   a          
          !   �      �     �   >      �     �   /   L      a         	                n  D            n  �            !  �   #      !  �   #   .        #   i      �      �   #   �   !   �   !   �   !   i   a           �         �      �     �   /   A                     #  �   !  �            #  �   !  �            #  �   !  �                     b                  n        ��c�Y\�9��'�         !  �   #      !  �   #   .        #   i   !   �   !   �   !   i   a           �         �      �     �   /   A                     #  �   !  �            #  �   !  �            #  �   !  �                     b         !   �      �   W      (   g            n  p            !  �   #      !  �   #   .        !   �      =   ����       W      (   g            n  �            !  �   #      !  �   #   .   !   �      �     �   a          �`��h�
�㜁8   
          !   �   !        �     �   /   L      a         	                n  8            !  �   #      !  �   #   .         !   �   )   6             !   �   )   6               �   )   6   0            �   )   6   `         !   �   )   6   p         !   �   )   6   �   !   3   !     a           �         �      �   A                     #  �   !  �            #  �   !  �                     b                  6                6         �P�wo��d9A�         6                6   0            6   @            6   P            6   `            6   p            6   �      x      
      #  �   !  �      	      #  �   !  �      	      #  �   !  �      	      #  �   !  �      	      #  �   !  �      	      #  �   !  �      	      #  �   !  �      	      #  �   !  �      	      #  �   !  �      	         
   	   b   y   	            n  d            !  �   #      !  �   #   .   !   �      �   ���$����' ��     �   a          
          !   �   !   �     �   >      �     �   /   L      a         	                 n  �      !      !  �   #      !  �   #   .   !   ,      �      �   a   /      
       !   �      �     �   /   L      a         	       !   -      �      �   a   /      
       !        �     �   /   L      a         	          ,      -      M      L         �   I   #   �      �      �         #   n  ,      $      !  �   #      !  �   #   .   !   �j����j	u+g   �      �     �   a          
          !   �   !   �     �   >      �     �   /   L      a         	          %      n  �      &      !  �   #      !  �   #   .   "   1      !   �      �     �   /   a         	       "   1      !   �      �     �   /   a         	                       (         (   >        (   $              (   �             2            #  �   !  �            b         !   �   "   1         �     �   /   a         	       ���������   !   �   "   1         �     �   /   a         	          '      n  X      "         #      n  �      (      !  �   #      !  �   #   .   !   �      �     �   a          
          !   �   !   �     �   >      �     �   /   L      a         	          )      n  L      *      !  �   #      !  �   #   .   !   ,      �      �   a   /      
       !   �      �     �   /   L      a         	       !   -      �      �   a   /      
       !         �     �   �,w���   /   L      a         	          ,      -      M      L         �   I   #   �      �      �         ,      -      !  �   #      !  �   #   .                   (         (   >     !   (   $           "   (   �             2            #  �   !  �            b            .         +         ,      n  �      /      !  �   #      !  �   #   .      �      �   =      	         #      M      L         �   I   #   �      �      �         1      2   ��K���YC�4�      !  �   #      !  �   #   .   !   �      �     �   a          
          !   �   !  $      �     �   /   L      a         	          3         4      1         0      n   l      5      !  �   #      !  �   #   .      �      �   =      	         %      M      L         �   I   #   �      �      �         7      8      !  �   #      !  �   #   .   !   �      �     �   a          
          !   �   !  &      �     �   /   L      a         	          ��V�l@�b�ǒ�   9         6         7         4      n  !4      :      !  �   #      !  �   #   .   "   1         �      �     �   /   a         	       "   1      !   �      �     �   /   a         	       "   1   #   !   �      �     �   /   a         	       "   1   2   !   �      �     �   /   a         	       "   1   =   !   �      �     �   /   a         	                       (         (   >     '   (   $           (   (   �             2            #  �   �ҧ���@�Gv�o�   !  �            b            �   "   1         �     �   /   a         	       !   �   "   1         �     �   /   a         	       !   �   "   1   #      �     �   /   a         	       !   �   "   1   2      �     �   /   a         	       !   �   "   1   =      �     �   /   a         	          ;      n  #�      <      !  �   #      !  �   #   .   !   ,      �      �   a   /      
          �      �     �   /   L      a         	       !   -      �   ����>w�Ē      �   a   /      
       !  )      �     �   /   L      a         	          ,      -      M      L         �   I   #   �      �      �         >      ?      !  �   #      !  �   #   .                   (         (   >     *   (   $           +   (   �             2            #  �   !  �            b            @         =         >      n  %�      A      !  �   #      !  �   #   .   !   ,      �      �   a   /      
          �      �      �.�q����;4l  �   /   L      a         	       !   -      �      �   a   /      
       !  ,      �     �   /   L      a         	          ,      -      M      L         �   I   #   �      �      �         C      D      !  �   #      !  �   #   .            �   )   6       !   3   !  -   a           �         �      �   A                     #  �   !  �            #  �   !  �                     b                  6          x            #  �   !  �      ����k�7�e         b   y         E         B         C      n  &�      F      !  �   #      !  �   #   .   !   �      �     �   a          
          !   �   !  .      �     �   /   L      a         	          G      n  '      H      !  �   #      !  �   #   .     /   =   ����       #   �      I         �      n  't   n  '�      J      !  �   #      !  �   #   .      �   =      	         0   <              #   �      �   =   ����       #   �      K      n  (<      �1C��p���Y�   L      !  �   #      !  �   #   .      �   =              W        �   N      4   #   �         !  3   !  2   !   �   !  1   c   w                    !   ,      �      �   a   /      
          �      �   >      �     �   /   L      a         	       !   -      �      �   a   /      
       !  4      �     �   /   L      a         	          ,      -      M      L         �   I   #   �      �      �         N      �      M         N      n  )      O   �J�������k��      !  �   #      !  �   #   .      �   =              W        �   N      4   #   �         !  7   !  6   !   �   !  5   c   w                    !   ,      �      �   a   /      
          �      �   >      �     �   /   L      a         	       !   -      �      �   a   /      
       !  8      �     �   /   L      a         	          ,      -      M      L         �   I   #   �      �      �         Q      �      P         Q      n  )�      R      ��:�!"��n'H   !  �   #      !  �   #   .   !   �         �   L      N        �   a          
             �     �   /                �      L      a         	       >   #   �      T         �     �   ?      #   �      0      �   L         L         U       U      �   !   �         T      V      U         �     �   >   #   �      V         �      !   �   @   K      #   �      �     �   /   !  9     �   >      L      a         	          �      �     �   a       ��,J��[���g      
             �   !   �      �     �   /   L      a         	          S         �      n  *0   n  *�      W      !  �   #      !  �   #   .   !   �         �   L      N        �   a          
             �     �   /                �      L      a         	       >   #   �      Y         �     �   ?      #   �      0      �   L         L         Z       Z      �   !   �         Y      [      Z         �     �   >   #   �      [         �      ����i���|��}\   !   �   @   K      #   �      �     �   /   !   �     �   >      L      a         	       !   �      �     �   a          
          !   �   !   �      �     �   /   L      a         	          X      n  *�      \      !  �   #      !  �   #   .           �   >         �   N        �   a          
                �     �   /   (   �   !   �         !  :   )   �       !   �         !  ;   )   �   0         �     �   /   )   �      c   �             !   �03�Z�t���   �      �     �   /   >      (   g      ]      n  +�      ^      !  �   #      !  �   #   .   !   �     �   >      g   V   
   #   �      �   =      	         <      M      L         �   I   #   �      �      �         `      a      !  �   #      !  �   #   .                   (         (   >     =   (   $           >   (   �             2            #  �   !  �            b            b         _         `      n  .|      c      !  �   #      ��BI>�D&��T   !      #   .   !   ,      �      �   a   /      
          �      �        /   L      a         	       !   -      �      �   a   /      
       !  ?      �     �   /   L      a         	          ,      -      M      L         �   I   #   �      �      �         e      f      !     #      !     #   .                   (         (   >     @   (   $           A   (   �             2            #  �   !  �            b            g         d   �YTt*�t0�c�/�         e      n  0      h      !     #      !     #   .   !   ,      �      �   a   /      
          �      �        /   L      a         	       !   -      �      �   a   /      
       !  B      �     �   /   L      a         	          ,      -      M      L         �   I   #   �      �      �         j      k      !     #      !     #   .      �      �        a          
             �      �      �     �   /   L      a         	          ��p���T�[��5   l         i         j      n  2d      m      !     #      !  	   #   .   !   �      �     �   a          
          !   �   !   �     
   >      �     �   /   L      a         	          n      n  2�      o      !     #      !     #   .   !   �      �     �   a          
          !   �   !   �        >      �     �   /   L      a         	          p      n  3�      q      !     #      !     #   .   !   �      �     �   a          
          !   �U7vu����.��n   �   !  C      �     �   /   L      a         	          r      n  3�      s      !     #      !     #   .   "   1      !   �      �     �   /   a         	                       (         (   >     D   (   $           E   (   �             2            #  �   !  �            b         !   �   "   1         �     �   /   a         	          t      n  4X      u      !     #      !     #   .   !   �         �   L      N        �   a          ������d�,��   
             �     �   /             !  F      L      a         	       >      �     �   /   !   �     �   >      L      a         	       !   �      �     �   a          
          !   �   !   �      �     �   /   L      a         	          v      n  4�      w      !     #      !     #   .   j   �   l����       j   �   l����       "   1      !   �      �     �   /   a         	                       (         (   >     G   (   $           H   (   ��Es�n���9   �             2            #  �   !  �            b         !   �   "   1         �     �   /   a         	          x      n  5    k   �   l����       k   �   l����          y      �         z     	         z   !   z     	      	   c   {                 z         {      !     #      !     #   .   "   1      !   �      �     �   /   a         	                       (         (   >     I   (   $           J   (   �             2            #   �*���kPcbPn�  �   !  �            b         !   �   "   1         �     �   /   a         	          |         y   n  5�      �         z     	         }   !   z     	      	   c   {                 }         ~      !     #      !     #   .                   (         (   >     K   (   $           L   (   �             2            #  �   !  �            b                     y      n  7x      �      !     #      !     #   .   !   �      �     �   ����F7�wy�-   a          
          !   �   !  M      �     �   /   L      a         	          �      n  7�      �      !     #      !     #   .   "   1         �      �     �   /   a         	       "   1      !   �      �     �   /   a         	       "   1   #   !   �      �     �   /   a         	       "   1   2   !   �      �     �   /   a         	       "   1   =   !   �      �     �   /   a         	       "   1   H   !   �      �     �   /   a         	       ���T�8�|���o                   (         (   >     N   (   $           O   (   �             2            #  �   !  �            b            �   "   1         �     �   /   a         	       !   �   "   1         �     �   /   a         	       !   �   "   1   #      �     �   /   a         	       !   �   "   1   2      �     �   /   a         	       !   �   "   1   =      �     �   /   a         	       !   �   "   1   H      �     �   /   a         	          ���'֑��z��   �      n  :�      �      !     #      !     #   .   !   �         �   L      N        �   a          
             �     �   /                �      L      a         	       >   #   �      �         �     �   ?      #   �      0      �   L         L         �       �      �   !   �         �      �      �         �     �   >   #   �      �         �      !   �   @   K      #   �      �        /      �     �   >      L      a         	          ��d��C-��N�5�   �        N      /   #   �   !   �         �   L      N            a          
             �             !   �      M      a         	       >   #   �      �         �     �   ?      #   �      0      �   L         L         �       �      �   !   �         �      �      �         �     �   >   #   �      �         �      !   �   @   K      #   �      �     �   /   !  P     �   >      L      a         	       !   �      �     �   a          
       ���)e����      !   �   !   �      �     �   /   L      a         	          �      n  ;`      �      !  !   #      !  "   #   .            �   )   6             !   �   )   6            !   �   )   6             !   �   )   6   0         !   �   )   6   @            �   )   6   P            �   )   6   `            �   )   6   p            �   )   6   �            �   )   6   �            �   )   6   �            �   )   6   �            �   )   6   �            �   ��r.�OM��j   )   6   �            �   )   6   �   !   3   !  Q   a           �         #      �   A                     #  �   !  �            #  �   !  �                     b                  6                6               6                6   0            6   @            6   P            6   `            6   p            6   �            6   �            6   �            6   �            6   �            6   �            6   �      x      �d�xBfF.Q�5G         #  �   !  �            #  �   !  �            #  �   !  �            #  �   !  �            #  �   !  �            #  �   !  �            #  �   !  �            #  �   !  �            #  �   !  �            #  $   !  $            #  %   !  %            #  &   !  &            #  '   !  '            #  (   !  (            #  )   !  )                     b   y         �      n  >�      �      !  *   #      !  +   #   �*~��QvgPxh   .   "   1      !   �      �     �   /   a         	                       (         (   >     R   (   $           S   (   �             2            #  �   !  �            b         !   �   "   1         �     �   /   a         	          �      n  ?H      �      !  ,   #      !  -   #   .                   (         (   >     T   (   $           U   (   �             2            #  �   !  �            b            �      n  @      �  �t���-:�      !  .   #      !  /   #   .   !   �         �   L      N        0   a          
             �     �   /             !  V      L      a         	       >   #   �      �         �     �   ?      #   �      0      �   L         L         �       �      �   !   �         �      �      �         �     �   >   #   �      �         �      !   �   @   K        �   N      /   #   �     �   >      �     �   /      �     �   >      L      a         	  βyq]���M�҇          �     �   N      /   #   �   !   �         �   L      N        1   a          
             �             !   �      M      a         	       >   #   �      �         �     �   ?      #   �      0      �   L         L         �       �      �   !   �         �      �      �         �     �   >   #   �      �         �      !   �   @   K        �   N      /   #   �     �   >      �     2   /   !  W     �   >      L      a         	         �,[5e�����   �     2   N      /   #   �   !   �         �   L      N        3   a          
             �             !   �      M      a         	       >   #   �      �         �     �   ?      #   �      0      �   L         L         �       �      �   !   �         �      �      �         �     �   >   #   �      �         �      !   �   @   K        �   N      /   #   �     �   >      �     �   /      �     �   >      L      a         	          �     �\�����|�<$.  �   N      /   #   �   !   �         �   L      N        4   a          
             �             !   �      M      a         	       >   #   �      �         �     �   ?      #   �      0      �   L         L         �       �      �   !   �         �      �      �         �     �   >   #   �      �         �      !   �   @   K      #   �      �        /      �     �   >      L      a         	          �        N      /   #   �   !   �        �
'�Z� �e���   �   L      N        5   a          
             �             !   �      M      a         	       >   #   �      �         �     �   ?      #   �      0      �   L         L         �       �      �   !   �         �      �      �         �     �   >   #   �      �         �      !   �   @   K      #   �      �     �   /   !  X     �   >      L      a         	       "   1      !   �      �     5   /   a         	                       (        ]7��ۇ���j��   (   >     Y   (   $           Z   (   �             2            #  �   !  �            b            �      n  A�     [   #   "            �      n  C0   n  C�      �      !  6   #      !  7   #   .      �      �         �      �      !  8   #      !  9   #   .                   (         (   >     \   (   $           ]   (   �             2            #  �   !  �            b            �         �         �      n  D�      �      !  x��#�v�p�  :   #      !  ;   #   .        #   �      �      n  E�      �      !  <   #      !  =   #   .   !   3   !  ^   a           �         >      �   A                     #  �   !  �            #  �   !  �                     b                  6                6               6                6   0            6   @            6   P            6   `      x            #  �   !  �            #  �   !  �            #  �   !  �           �{N��5��gz�   #  �   !  �            #  �   !  �            #  �   !  �            #  �   !  �                     b   y         �        _   #   "                                       .               n  G�      &   a           �         ?     l   A                     #  �   !  �            b            �      �         e      f   +   j  u   j  {   j     g   E      z     	            !   z     	      	   c   {                       !  	�i��ls&&�;   E      F          #   :   #   =   !   �                  �   L      N        @   a          
             E   )   �         �   )   �   0      �   )   �   A   a           �         A     m   A                     #  B   !  B            b         !   �      �   @      �   L        C   /   L               !   9      �   c   7                       !   �      �   @      �   L        D   /   L               !   <      �   c   7                      
�h�i<8����                     e   +   f      j  u   j  {   j     g   v      v      o          q      a           �         E      �     F   /   A                     #  G   !  G            b                           e          �                           �                                    7   +         6              w   L      {   Y      �   f      +   n             ~   �     �   �     �   �     �   �                      ��������@@@@@@@@@@@@@@  Г|�)�~���@@@@@@@@�                                                                                                                            |   ��                                                                       ��0                                                                                                                                                                                                                                                                       �                         �s��fJN(F��                                                "                              
               :                  $           @     �� ��                                                                                                                                                                                                                                                                                                                                                      ��R�=�'P<                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �s�Xo   !�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   !�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   "    � ���         ?�G7�  '*,	�        ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ��۪���&H�uP                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �s�Xo   "@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   "`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   "�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   "�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   "�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   "�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   #  �����                                  0                                      P  `  P ���������� @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                ��������@@�����@@@@@�����@@@@@@@@@@@@@@@@            \���@@@@@@@@@@@@@@@@\������@@@��      �          @@@@@@@@@@@@@@@@@@@@@�@@@@@@@@@@@@@@@��������������������������������������������@@@@��������@@�������@@@@@@@@@@@@@@@@@@                                @@                      �       �          ������@@@@����@@@@@@          ����G���=��'L�  �y�OmX&���������@@@@����@@@@@@          ������@@@@@@@@@@������@@@@����@@@@@@          D�����9{���.���������@@����@@@@@@          ��������@@@@@@@@                                                                                                                                                                                                                                                                                                                                                                                  �o�S�5��O�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �s�Xo   #`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   #�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   #�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   #�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   #�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo   $    `� ���         ��  �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           !�*�n]1�&:4 8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "�s�Xo   $@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   #�s�Xo   $`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   $�s�Xo   $�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   %�s�Xo   $�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   &�s�Xo   $�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   '�s�Xo   $�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   (�s�Xo   %                                  ���@⨔���@あ��       *  �   @  `  
@   T  �  �            ���� ��������@@                     P������ P�������� P������ P���� P������� P������� P���� P������� P� P��� P������� P������ P���������� P������ P������ P����� P���� P������ P������ P���������� P�������� P��������� P��� P������� P������� P��������� P������ P������ P������ P������� P�������� P������ P���� P������ P��������� P������� P���� P���������                           �                       ����          )�Y�i��� �\                                 ����                  0                      ����                  `                       ����                  �   @                                        �                                            �     �            
   ����                                                              P            �                            �   �   �      �                            �              �                            �                   *�/^�j�%�~�Ux                           P   P      �    
                        @                         	                  p   P   P      �          
                  �   0   0      �                            �                                             �   �      �                            0   P   P      �                            `   0   0      �                            �                                         �   P   P      �                            �  �  +Ir�B#��ߔ  �      �                                8   8      �                            P            �                            �   P   P      �                            �              �                            �                                            x   x      �                            @                                         p            �                            �   �   �      �                            �  0  0      �                    ,������oW�                                                    0              �                            `              �                            �              �                             �   H   H      �          !                  �  @   @       �          "                  	                         #                  	P            �          $                  	�            �          %                  	�                       &                  	�  (  (      �      -�{-��Bլ�      '                  
   P   P      �          (                                           E                  
�  
�   0  �       E                 
�  
�     �                                               �   E                                 �  �   �   �          
                 0  �  p   �   �                           `  �  �   ~   �                           �  �  P   l   �                                       d   �                                   .�x+��$&�{1�  �   v   �                              P     �   �                                   �   �   �          	                         @   �   �                           �  @  0   �   �                           �    �   �   �                                   �   �   �                                       �   �                           p  �  �   �   �                                   `   �   �                                   �   �   �                   /����S̽��Fh             P  p     �                           0  �  �   �   �                           `  �  P   �   �                                       �   �                                   �   �   �                           �          �                                   �     �                                   @     �          "                 �  �  �  e   �                           �  @  0  B   �                           �    �  /   �      0�-h�[���3.�                               �  &   �                                      :   �                            p  �  �  R   �                                   `  J   �          !                         �  [   �          &                    �  	�  �   �          $                 0  `  	P  s   �          #                         	   m   �          %                         	�  {   �          '                     �  	�  �   �          (                         1B/�mw��r��  
  �   �       e                              �                                                                                                                                                                                                                                                                                                                                                                                                       E  �              
�               e                              d  2�p�?�9��8�              �  �  0                              �      X  �              |  �      \      �          x            ,          t      �      �                                  P                  �  `                              4      �                                          �  �          �                      �  �                      T           �  x              
�               �  �                              ~  �              0               l  �          3	q�i0� ]r�H      `               d                �               v  ,              �               �  P              �               �  t                              �  �              P               �  �              �               �  �              �               �                �               �  (                             �  L  �          @               �  p              p               �  �              �                �              �               �  �                 4�[�O�B���j5�               �                 0               �  $              `               �  H              �                l              �                �              �                �  <                         e  �              P              B  �              �              /     �          �              &  D              �              :  h  8                        R  �              @              J  �              p              [  �              �          5�r�iF��K1�O�      �  �              �              s    �                         m  @  �          0              {  d              `              �  �              �              �  �              �                    ���@�� �$                   ����@�����@����@  ��     �`               @  �`  �   �@  �`    �@����  � \����@@@@@@@@@@@@@@@@@@@@@@@@@\����@@@@@@@@@@@@@@@@@@@@@@@@@\��@@@@@@@����`�@@@@@@@@@@@@@@     %�������������   ����                                            �����@������@@@@  6��e�d��N��      0          @����nnnnnnnn����@����������@P��   �          �  �`��@Ӊ�����@剅�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\�   %@    ������������� �H��������  �   �������������@����@@@��@  �@     �  � ����@�������@������@@������@@@@@@@@@@@@@@@@@@Ö�����@Ӂ������@@@@@@@@@�������a��������@@@@@@��������@��a��a��@��z��z��@@@@@@@@@ׁ��@@@@� @י�����@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@z@@@��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@Ӊ�����@K@K  7n,Wӳ�,����@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@z@@@@@�������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @▤���@����@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@z@@@������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@Ӊ�����@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@z@@@@@�������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @▤���@������@����@@K@K@K@K@K@K@K@K@K@K@K@K@K@z@@@��������@@@��a��a��@��z��z��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  8�(���-i��R@@@@@ @▤���@��������@�������@K@K@K@K@K@K@K@K@K@K@K@z@@@\����@@\��������@@\��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @䢅�@�������@@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@z@@@\�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @י�����@�������@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@z@@@\���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @ą�����@����������@�����@@K@K@K@K@K@K@K@K@K@K@z@@@\��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  9��8��o@�2B@@@@@@@@@@@@@@@@@@@@@@@@@ @����������@�����@@K@K@K@K@K@K@K@K@K@K@K@K@K@K@z@@@\������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @م�����@�������@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@z@@@\��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @す���@�������@@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@z@@@������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @���������@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@z@@@\���������@@@@@@@@@@@@@@@@@@@@@@@@@@  :7��f�U�H4��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @▙�@��������@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@z@@@\���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @Ӂ������@����������@K@K@K@K@K@K@K@K@K@K@K@K@K@z@@@\������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @ㅧ�@@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@z@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @֗����������@@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@z@@@\����@@@@@@@@@@@  ;�:�x�e`-q�a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @ą�������@����@@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@z@@@\����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @ŕ����@�����������@����������@K@K@K@K@K@K@K@K@z@@@\���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @⣖����@�����@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@z@@@\������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @Ö������@@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@K@  <�2�n"s�2Jz@@@���@�⅙���@Ö�����@Ӂ������@Ö������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@Ö�����@Ӂ������@▤���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @������@@\KKKNKKK@�@KKKNKKK@�@KKKNKKK@�@KKKNKKK@�@KKKNKKK@�@KKKNKKK@�@KKKNKKK@�@KKKNKKK@�@KKKNKKK@�@KKKNK@@����@@@@@@@@@@@@@@@@@@@@@ @@@@���`@@@@@@@@@@@@@@���@@@@@@@@����MP����@P���@P������@P�������@P�������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@@���@@@@@@@@@@@@@@@@@@@@  =��3�6�
�r� i@@@@@@@@P��������@P��������@P���������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@P����������@P���������@P���������@P����@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@P����������@P���������@P������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@@���`@@@@@@@@@@@@@@���������@@����M}ǉ������@Ö���������@����@`@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@@���  >�q�L�ru�I�@@@@@@@@@@@@@@@@@@@@@@@@@@@@����������|�����K��}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@@���`@@@@@@@@@@@@@@���@@@@@@@@���MP����]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@@���`@@@@@@@@@@@@@@���@@@@@@@@���MP���]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@@���`@@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\���]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@  ?kjy��CE�X�@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP�������]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP�������]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP��������]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP��������]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  @˫=����zSq��@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP���������]@����M\���]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP����������]@����M\���]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP���������]@����M\���]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP���������]@����M\���]@���M�]@@@@@@@@@@@@@@  AWb^pH�Yk�v@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP����]@����M\���]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP����������]@����M\���]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP���������]@����M\���]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@��  BG����IX��J���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP�������]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP����]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP��  Cl�&^rdMw�E������]@����M\����]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP�������]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@  D��R�'����@@���@@@@@@@@���MP������]@����M\����]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP��������]@����M\����]@���M����]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@���M���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@   EP���D��Klӑ�@@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP����]@����M\����]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP�]@����M\���]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP�������]@����M\����]@���M���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP���]@����M\����]@���M���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a�  F�[�^sl>d3�?��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP����]@����M\����]@���M�]@�����M�}��}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@���M���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP�������]@����M\����]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@  G7"��ޗYʺ�P@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP����]@����M\����]@���M���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP�����]@����M\����]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@���M��]@@@@@@@@  H!��Or�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���@@@@@@@@���MP�������]@����M\���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@������@@@@@�����M�������]@����M����@������M�����]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@����`@a\@ǅ�@���@����������@��@���@�������@����@@@  I_����B�����@@@@@@@@@@@@@@@@@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@����`@a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@������@@@@@���MP����]@�����M}�}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@��@@@@@@@@@����MP���@~@}\}]@����M�������@���MP�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����@@@@@@@@@@@@@@@@@@@@@@@@@@  J����m�eb�D@@����MP����]@���MP������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@����@@@@@@@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@������@@@@@���MP�������]@�����Ml���MP���@�@��]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@������@@@@@���MP����]@�����Ml���MP���@��@��]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@  K!��CQE�Ǵ@@@@@@@@@������@@@@@���MP������]@�����Ml���MP���@��@�]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@������@@@@@���MP�������]@�����MP������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@������@@@@@���Ml���MP������]]@�����MP�������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@  LFTs�I ��{�ٝ@@@@@@ @@@����`@@@@@@@@@@@@@@������@@@@@���Ml���MP������]]@�����M����]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@������@@@@@���MP������]@�����M�}����������������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@����@@@@@@@���M��������]@����MP��������@P������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@}��������}@P���@}@}@}@}@P����@P������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  M�Aӣ>����a��a��@@@@@@@@@@@@@@@@@@ @@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@P������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@������@@@@@���MP�����]@�����Ml���MP������@�@�]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@��@@@@@@@@@����MP�����@\��@}@}]@����M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@������@@@@@���MP������]@�����Ml���MP������@��@��]]@@@@@@@@@@@@@@  N8��=b��H%�~�@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@���������@@�����MP�����]@����M�������]@������MP������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������M\������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@a\```````````````````````````````````````````````````````  O6�Ӕ��=���5`````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@����`@a\@È���@���@������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@����`@a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@������@@@@@���MP�������]@�����Ml���MP��������@���@��]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@��@@@@@@@@@����MP�������  Pb���fTS�����@\��@}\���}]@����M���������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@�����M�������]@����M�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@������M}◖��@��@���@\���}]@�������M\������]]@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@����`@a\@È���@��@���@�  QN;B�n��ԋy{��������@��@����������@��@���@�����@@@@@@@@@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@����`@a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@��@@@@@@@@@����MP������@~@`�]@����M������@���MP�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@�����M\����]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@���  R �����7-A�`@@@@@@@@@@@@@@����@@@@@@@���M��@����MP������@~@�]@����M������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@���MP�������]@�����M\����]]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@��������@@@����MP����]@���MP������aP����aP�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@������MP�������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@  Sv��U��s��1@@@@@@@@@@@@@ @@@����`@a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@����`@a\@È���@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@����`@a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@����`@a\@ׁ��@�������@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  T�9�tЕ�j��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@��@@@@@@@@@����MP�������@~@}@}]@����M���������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@�����M�������]@����M�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@������M}ׁ�������@�������@�������}]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������M\������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@  U���ؾ�#�ǋ��@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@a\@ą�����@����@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@��@@@@@@@@@����MP�������@~@}\������}]@����M����@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@���M��������]@����MP�������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@����`@a\@È���@ׁ��@���������@\a@@@@@@@@@@@@@@@@@@@@@@@@  VM�Z�10zsǪ�,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@����`@@@@@@@@@@@@@@������@@@@@���MP����]@�����M}�}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@������@@@@@���MP�]@�����M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@��������z@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@������@@@@@���MP�  W`�SJQ���*�]@�����MP�@`@�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@��@@@@@@@@@����Ml���MP�������@P�@�]@~@}a}]@����M����@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@������M���������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@��@@@@@@@@@����Ml���MP�������@P�@�]@~@}@}]@����M����@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@  X���Z���!#r�@@@@@@@@@@@@@@@@������M��������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@������@@@@@���MP�������]@�����MP�������@\����@}a}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@���������z@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@������@@@@@���MP�������]@�����MP�������@\����@P����]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@  Y�Ѽ	)ݎC��� @@�����`@@@@@@@@@@@@@@�������@@@@���M}����}]@����MMP�������]@MP������]]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@������Ml���MP������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@��@@@@@@@@@����Ml���MP������]@\��@�]@����M���������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@�����M�������]@����M�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a  Z[4ٻ/�NE�����@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@������M}晖��@ׁ��}]@�������M\������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@a\@È���@���@Ձ��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@  [�'�eW�p��B@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@a\@�������@�������@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@��@@@@@@@@@����MP�������@~@}@}]@����M���������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@�����M�������]@����M�������]@������M}���@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@����@�������}]@�������M\������]]@@@@@  \:�����|�u9�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@a\@ą�����@�������@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@��@@@@@@@@@����MP�������@~@}\����}]@����M������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@���MP�������]@�����MP����]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@a\`````````````````````````````````````````  ]�w��+�p�S```````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@a\@Ö��@���@◖��@����@�@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@a\@ǅ�@���@�����@����@����@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@������@@@@  ^w��'Z�+O.�@���MP������]@�����Ml���MP��������@���@�]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@������@@@@@���MP������]@�����Ml���MP��������@���@�]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@a\@���@�@������@���@����@�����@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@������@@@@@���MP����]@�����M}�}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@@@@  _$�����.p��G@@@@@@@@@@���������@@������M�����]@������MP�������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@������@@@@@���MP������]@�����M}�}@\���@P�������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@������@@@@@����M����a��������]@���MP������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@������@@@@@�����M�������]@����M������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@  `� ���B<�z@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@����M����a��������]@���MP������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@������@@@@@�����M�������]@����M���������@�����M�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@����M�������]@������M}���@����@���@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@�����}]@�������M\������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  a�}z���[��aj@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@a\@Ö��@���@���������@����@���@������@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@������@@@@@���MP����]@�����M}�}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@�������@@@@����MP����]@������M����a��������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@���MP������aP����aP�������]@N@@@@@@@@@@@@@@@@@@@@@  b���|V�j�@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@������MP�������]@�����MP������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@������M\���]@�������M\����]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@a\@Ù����@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  cO��x%�gtΩ|�@@@@@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@������@@@@@���MP���]@�����MP�������@\����@P�������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@\����@}K���}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@����@@@@@@@���M��������  dΆ͋k�e���O]@����MP����@P������@P������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@P������@P���@P��������@P��������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@P���������@P����������@P���������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@P���������@P����@P����������@P���������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@  e�=��ɖ1g�W@@@@@@@@@@P������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@a\@ㅙ������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@���  f��#b(�՚0�<��`@a\@م����@���@���������@����@��@���@�����@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@����@@@@@@@����M����a��������]@���MP������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@������@@@@@����M\����]@�����M\���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@a\@⅕�@�@����������@�������@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  g=w���� ���@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@���������@@�����M�������]@����M�������]@������M}◖��@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@����}@\����@P����@\����@}���������@����}@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@\����@P�������@\����@P�������@\����@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@}K���}]@�������M\����]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  h���*��J�Bh@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@a\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@a\@ř����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@a\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\  ir6���O���a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@�����z@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@��@@@@@@@@@����MP�������]@����M���������@�����M�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@����M�������]@�������M\������]]@a\@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@��������@�����@@@@@@@@@  j�K��m���.�@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@������@@@@@���MP�������]@�����M}�}]@a\@���@������@��@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@�����@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@����@@@@@@@���M��������]@����M}@@@@}@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@�}�  k�OEY0S�N?�����������������������������}@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@�}�����������������������������������������N@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������������������������������������N@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@������������}@�}��������}@��������@\@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����@@@@@@@@@@@  lr5�
&%�p��@@@@@@@@@@@@@@@@@�}��������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@�����`@@@@@@@@@@@@@@������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��a��a��@@@@@@@@@@@@@@@@@@ @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\@\@\@\@\@@@�@�@�@@@�@�@@@�@�@�@�@�@�@@@\@\@\@\@\@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@Ù���@م�������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  m�P�^������@ @ą������@偙������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @Ձ��@@@@@@@@@@@@@@@@@@@@@@@@ą�����@@@@@㨗�@@@@@@@@@@@@Ӆ����@@@@@@م��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P������@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@���@@@@@@@@@@����@@@����@@@����@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P��������@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@@��@@@@@@@@@@@���@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@  nR�V�y�2�+�`@@@@@@@@@@@@@@@@@@@@@ @P������@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@@@�@@@@@@@@@@����@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P����@@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\���@@@@@@@@@@@@@@@@�@�@@@@@@@@@���@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P�������@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@@��@@@@@@@@@@����@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P�������@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\���@@@@@@@@@@@@@@@@�@@@@@@@@@�����@@�����@@@@@@@@  o;���6[V=�B�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P����@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@\����@@@@@@@@@@@@@@��@@@@@@@@@@@���@@@����@@@����@@�����@@�����@@�����@@�����@@@@@@@@@@@@@@ @P�������@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@@@�@@@@@@@@@@����@@@����@@@����@@@����@@@����@@�����@@@@@@@@@@@@@@@@@@@@@ @P�@@@@@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\���@@@@@@@@@@@@@@@@�@�@@@@@@@�����@@�����@@�����@@�����@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P���@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@\����@@@@@@@@@@@@@@��@@@@@@@@@  p��et�x`I�@@���@@@����@@@����@@@����@@@����@@@����@@@@@@@@@@@@@@@@@@@@@ @P�������@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@@��@@@@@@@@@@����@@@����@@@����@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P������@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@@@�@@@@@@@@@@����@@@����@@@����@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P����������@@@@@@@@@@@@@@@@@@@����@@@@@@\���@@@@@@@@@@@@@@@@�@�@@@@@@@@@���@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P������@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@  q,���{�'��@@@@@@@@@��@@@@@@@@@�����@@�����@@�����@@�����@@�����@@�����@@@@@@@@@@@@@@@@@@@@@ @P������@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@@��@@@@@@@@@@����@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P�����@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@@@�@@@@@@@@@@����@@@����@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P����@@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@@@�@@@@@@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P������@@@@@@@@@@@@@@@@@@@@@@@  r�D�H!e<�:�����@@@@@@\����@@@@@@@@@@@@@@��@@@@@@@@@@@���@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P������@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@@@�@@@@@@@@@�����@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P����������@@@@@@@@@@@@@@@@@@@����@@@@@@\���@@@@@@@@@@@@@@@@�@�@@@@@@@@@���@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P��������@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@@��@@@@@@@@@@@���@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P���������  s��nVa3�s�@@@@@@@@@@@@@@@@@@@@����@@@@@@\���@@@@@@@@@@@@@@@@�@�@@@@@@@@@���@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P���@@@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@���@@@@@@@@@�����@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P�������@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@@��@@@@@@@@@@@���@@�����@@�����@@�����@@�����@@�����@@@@@@@@@@@@@@@@@@@@@ @P�������@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@@��@@@@@@@@@@@���@@@����@@@����@@@����@@�����@@�����@@�����@@����  t�b{��1َ���/�@@����� @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�����@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P���������@@@@@@@@@@@@@@@@@@@@����@@@@@@\���@@@@@@@@@@@@@@@@�@�@@@@@@@@@���@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P����@@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ \@�������@��@@偙�����@P����@��������@���@���@��������@��K@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  u8j]�!*�^^�@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P������@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@@@�@@@@@@@@@�����@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P������@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@@@�@@@@@@@@@@����@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P������@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@@@�@@@@@@@@@�����@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P�������@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@@@�@@@@@@@@@�����@@�����@  v��Y�qO7t>@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P��������@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@����@@@@@@@@@@����@@@����@@�����@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P������@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@\���@@@@@@@@@@@@@@@@�@�@@@@@@@@@���@@@����@@@����@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P����@@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@@@�@@@@@@@@@@����@@@����@@�����@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P������@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@���@@  w��Z42S��@@@@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P���������@@@@@@@@@@@@@@@@@@@@����@@@@@@\���@@@@@@@@@@@@@@@@�@�@@@@@@@@@���@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P�������@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@���@@@@@@@@@�����@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P����@@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@\����@@@@@@@@@@@@@@��@@@@@@@@@@����@@@����@@@����@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @P���������@@@@@@@@@@@@@@@@@@@@����@@@@@@\��  x?S뺃�!L�)�@@@@@@@@@@@@@@@@�@�@@@@@@@@@���@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @ą�����@Ӂ����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @Ӂ���@@@@@@@@@@@@ą�����@@@@@م��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @���������@@@@@@@@@�����@@@@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @�����@@@@@@@@@@@@@�����  y�8�����D@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @��������@@@@@@@@@@�����@@@@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@@@@@@@@@@@@@@@@@@@\@\@\@\@\@@@�@�@�@@@�@�@@@�@�@�@�@�@@@�@�@�@�@�@�@�@�@�@@@\@\@\@\@\@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\@\@\@\@\@@@�@�@�@@@�@�@@@�@�@�@�@�@�@�@�@�@�@�@@@\@\@\@\@\@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  nnn  z[ps1�6�e�����@����������@     @       �`����  @       �    �    �  &  �  0  �  :  �  D  �  	N  	�  
X  
�  b  �  l  �  v  �  �    �    �    �  #  �  -  �  7  �  A  �  K  �  U  �  _  �  i  �  s  �  }    �    �    �     �   *   �  !4  !�  ">  "�  #H  #�  $R  $�  %\  %�  &f  &�  'p  '�  (z  (�  )�  *	  *�  +  +�  ,  ,�  -'  -�  .1  .�  /;  /�  0E  0�  1O  1�  2Y  2�  3c  3�  4m  4�  5w  5�  6�  7  7�  8  8�  9  9�  :$  :�  ;.  ;�  <8  <�  =B  =�  {�A��JL�s  >L  >�  ?V  ?�  @`  @�  Aj  A�  Bt  B�  C~  D  D�  E  E�  F  F�  G!  G�  H+  H�  I5  I�  J?  J�  KI  K�  LS  L�  M]  M�  Ng  N�  Oq  O�  P{  Q   Q�  R
  R�  S  S�  T  T�  U(  U�  V2  V�  W<  W�  XF  X�  YP  Y�  ZZ  Z�  [d  [�  \n  \�  ]x  ]�  ^�  _  _�  `  `�  a  a�  b%  b�  c/  c�  d9  d�  eC  e�  fM  f�  gW  g�  ha  h�  ik  i�  ju  j�  k  l  l�  m  m�  n  n�  o"  o�  p,  p�  q6  q�  r@  r�  sJ  s�  tT  t�  u^  u�  vh  v�  wr  w�  x|  y  y�  z  z�  {  {�  |  |�  })  }�  ~3  ~�  =  �  �G  |�����鎩���  ��  �Q  ��  �[  ��  �e  ��  �o  ��  �y  ��  ��  �  ��  �  ������@����������@ �    �          � �������@⣁������@剅�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����`�@@@@@@@@@@@@@@\�   %@    <������������� k��������  � ������������@����������@ �      <     � ����  �` �       d        �        �        �        �                |        �        D        �                p        �        8   
     d        �        ,        �        X        �     }p�.
�q�^:5     L        �         l        !4        #�        %�        &�        '        't        '�        (<        )        )�        *0        *�        *�   
     +�        .|        0        2d        2�        3�        3�        4X        4�        5         5�        7x        7�        :�        ;`   
     >�        ?H        @        A�        C0        C�        D�        E�   
     G�   ���@����������@@      @        ~���La-�%  �@  �@@@@  �`����      nnnn���@����������@@         <     �`����@@@  @  �`        F      J      L      M      N      O      P      Q    	  R    
  S      T      U      X      Y      Z      [      ]      ^      b      e      j      l      n      v      y      {      |      }      ~      �      �       �    !  �    "  �    #  �    $  �    %  �    &  �    '  �    (  �    )  �    *  �    +  �    ,  �    -  �    .  �    /  �    0  �    1  �    2  �    3  �    4  �    5  �   ���s�rPx$�C�   6  �    7  �    8  �    9  �    :  �    ;  �    <nnnnnnnnnnnn���@�����@@@@@@@      X      ��������������  ����  �@     �`  �@      @������  ����                                                                                                                                                                                                                                                                                                                                                                          ���D��"{��o�  � ���         '*,	�  D               �  `                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ��yȼ*�&G� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��s�Xo   0@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   0`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   0�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   0�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   0�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   0�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   1                            0     p      0�����@����@�����\���������@@@@@@��������@@�����@@@@@            �������������   ��������        \���         �                \���     �  ��                                                                                                                  p           7�����@@@@@\����@@@@@          7����@@@@@@\����@@@@@          7��������@@\����@@@@@                                                                                                            ��ʜ���5��3                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��s�Xo   1@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   1`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   1�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   1�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   1�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   1�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   2  ������������@@@@@@@@@@@@@@@@@@@@@@                                   �   6 @ @                                                               �a�@������@����������@@@            ���� �s�TU�   �   �      �                                        ���V  �-X�s �                                                �-X�s �                                                                                                                                                                                          ���#O��`_��                                                                                                                                  @   @ #�R�*     0   0 '7nu     �   � C           ���V     p   p 쯉�           )^ʷ�           "                                                                                                                                                                                                                                                                                  ����\H�m.�	�b                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��s�Xo   2`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   2�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   2�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   2�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   2�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   3      � #�R�*   0     ���V  � ��������@@@@@@@@@@@@@@@@@@@@@@�       � @6 �s��JM� .�M��           
~6O   #�R�*       �s��S�                            �   �                               �                                       �              �ǁ ���        �                                                                                                                       ���� 0                                                                                                        ����t��LZWt,g                                                                                                                                   /ǉ������@Ö���������@����@`@����������|�����K��                   �#�R�* �       �#�R�*                                                             #�R�* @        #�R�* `#�R�*                 #�R�* �#�R�* �                                        #�R�* �                                                   �   X   `   �  �   �  �  �  �   �  �   �  p  `  P  @  ��2$�?���e�#�  0        �        #�R�* p������@@@@@@@@@@        #�R�* �D�����9{���.�        #�R�* ��������@@@@@@@@ P@�         ������@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@ P@�         ������@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@ P@�         ��������@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@�     �                                                     #�R�* �        #�R�* �#�R�* �                                #�R�* p   �   `        #�R�*   ���$���&i�              #�R�*      �        #�R�* @  `          #�R�* 	�  �  	@        #�R�* �     `                                                                                                                                        ������@@@@      \�@@@@@@@@                                                            @@@                                                                                                                                                                                        ��3�[T����C�                                                      @@@@@     ��������@@@@@@@@@@@@@@@@@@@@@@  \����@@@@@@@@@@@@@@@@@@@@@@@@@                                                                                                                                                                                                                                                                                                                                                                                               ��aM��`�׾V                                  @ ��                                         K                                      �a��������@@                                                                                                                                                                                                                  @@@                                                                                       @@                P  	   `  
0  p  �  �  P  �  p  �  �  	P     	`   p  ���I?�v��m�V8   p                   �         )�     �  P         '�     '    �         )      /P   �         )�   (                %m����m���m��������   $                      3                                                                                                                                                                                                                                                                                                                                              ��PV"�6�����}                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��s�Xo   4      �#�R�*  #�R�* �#�R�* �        #�R�* p#�R�* 0#�R�*   #�R�* 0#�R�* #�R�* �`  � �                 #�R�* p#�R�* �#�R�*                         � ߻Z                                        #�R�*  #�R�*  #�R�* 0#�R�* 8P#�R�* 6�                     �                                                                                                                                                                                                                                                  ��CS��F�fgH� `0000    000p`    �� 
 
����                                                                                                                                         �           #�R�*                                          '7nu                                          C                                                                                                                                                                                                                            �^�W�͆Ӛ�?H                                                                                                                                                                                                #�R�*                                                                                       �       �                                    �       �       �               �       �       �               �       �       �       �       �       �       �       �   '7nu      �       �       �       �       �       �     ��pO��|�%W�    �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �           #�R�* �             #�R�* �         �   #�R�* �             #�R�* �             #�R�* �         	    #�R�* �         
�   #�R�* �             #�R�* �         �   #�R�* �             #�R�* �             #�R�* �             #�R�* �             #�R�*           
    #�R�*          �   #�R�*         ��P�13���P�   :�   #�R�*          �   ����!���A��|�� (�!��`\  �A  < T� �!�3� `| �AڀSA݁��b h`}  �\  c^  �[P�;X�`��h�����_���?�����8`  8� K�`w  ����;@  ;  ; ��~��x;@��c�  K��`x  )  A�  �< x:����\ pb�  I�c"  N�!� � 0:�  �� @�^ @)� @� ��> 0� @~�@A� (�� @z�&�;>���Ȉ:�  ��  �� H  H�^ @;: {9  �� }9�@@� � �8H  {:$�*�� @z�&�;^�~���Ј� �� �> @;Y {Z  �^ @AՀ#K��h��z����`�;h�>�����^ 0�^�:��:���;5  ٨����z�' ꠁx(: 	|�z��b�  b�  �Y ;_��ꠁ{����{'   �g�!V�a���@�xz��(3 	|�zU�b�  c  �� "cC  c�  H  y�!  �����| �:_��;��� ����|�b�  c  � 28�  b�  bC  ~��bb  N�!A݁�Aڀc8!�� (|����N� !        ����#�R�* )��A���a�����|�� (�!�A`\  �A  < D� 3� �| �A݀�b h`}  �\  c^  �^j�^ ;@  �^h;@  �^��^ -  A� T�^ -� A���^ . @� ;@ �^�H  ��^ - @� ;@ �^�;@  �^�H |�^ -� A�,�^�.  A� \�
�{:�;  �  �< 0;��;^ �� (���{U' ꀁx(5 	|�z��b�  cU  �� "8�"�c  ~��c"  N�!;@ �^�:� ꠁ(|�b�  b�  �bH 
|�� /�����) @� l;@  �^�:� (  �G�/���(R�&� �(|�c6  b�  ��rH � @:���;^ � 8� �{W' ���x(7 	|�z��c6  cW  �� "b�  ~��c  N�!;@ �^�;  �> ���)� @� :�  ���:�  ���H 
<:�p; �ب�c  ; @@S9�{9 �8  �8 �8 �8 �8  �8 ":� �ר�b�  :�@@R����  ;U ڨ�cY  ; ��S��  � ���* @� :�  ���H  H  �� -  A� >�\�b���z��f��@b�@@���? \�c9��{9�g9��c9@@�>�;   � l;@ �^��m)� �@� (:�d���b�  :���R��z� ��  �� H  ;>d���c8  ;@��SZ�{Z �Y  �Y ���* �@� :�  ���H @:� ���� E) A�ԋm)� �A��;@ �^ EH ��>�.aA� ����  �G�$s����	�A-fA� ����z��� �x4�x�M�  A� \���z��� �{5�:� @���(|�b�  b�  � ���z��AՀ#� �| Hc4  � X�� ��  ��~��N� AՀ#�b| Hc:  � X�� �  ��~��N� ��֒� p��{:�� �������z��� �x9�x�N   A� ,���z��� �z��;; `���(|�b�  c5  �� :���b�  c�  H �AՀ#�b| Hc:  �� X� �  ��~��N� ��֒� p�< P;��;^ � H���{T' ���x(4 	|�z��b�  cS  �X ":�  �� 0�� 8c  ~��c"  N�!H  >�\�b���z��f��@b�@@����^m) �A�L>�\�b���z��f�@@b�@@���>`\�bs��zs�fs�@bs@@�~��
�z��;   �  ;   �>  ��f-4�W��|S�o:� ��P�^ �� ���^�:~���bt  :�@@R��z� ��  �� ;P:_�`;2 Pِ����{' �@�x(6 	|�{W�b�  c  �� �| `:_��:���\ X� �z�' ꠁx(7 	|�z��c  b�  �� "8� FbC  I�bb  N�!:� �Ȉ� z���� ��^
�zx��X  -� @� ;  �> pH  :�  �� p�� �*6  :� A� :�  -7  A� \��� b�A fzx�;@ @�X  ;8 ���c6  :�@@R��z� :� ~����  �� 	�� 	B ���� �� �� H 0:�  ��  :@  �_�p:~��@�zx' ���x(8 	|�z��cT  bu  �������p)���@� <�?�p�_��zx�~������V  *  A� ��p2� | H���pAՀ#K������� r�_��zy��! �� ������p  �7$�q�
����U)8 F@� ;@ F�_��H  ���p�����A vzv��! �����������z�  ��b�  c$  c  K�3�_������z��~r�Ӑ�bu  ���;  F�| H{  ��:� @bc  b�  b�  K�#;@  �^  :@ �^mAՀ#K��x>�\�b���z��f��@b�@@���AՀ#K���;?��c#  c�  H -AՀ#�^b| Hbt  � X�� ��  ��~��N� �^m)� �@� H  H  H  :� ����>�. @� ��~�- @� \�^ r-� �@� P� 0:���; �� (�@�{' � �x(5 	|�{:�cR  c  �W "8� �b�  ~��b�  N�!H  L� 0;?��; �\ (�`�{' ���x(2 	|�z�bv  c  �� "8�#)c#  I�b�  N�!H  T:�  ���^m* �@� ;  ��:` �~�  ��`�>�+J��a�H  :�  ���:�  ����>�:4Ȉ�
�z���R  H �; �`�{' ���x(7 	|�zӛbt  c  ��2;   �> Q;@ 1I�:[ x�؈:�p�����  ��  �� 	�� 	B ��;p:x����bu  :�@@R��z� ��  �� �� �� �� ;   �> D;@  �^ E:�  �� H:� �� P:@ �^ R;   � p:�  ��:�  ��:~�;3 \٘�c:  :�@@R��z� ��  �� :� f֘�b�  ; @@S�{ �  � :�ꀁ(|���r;[ ���(|�b�  cY  ��:{8�@�(|��^�:�  ������:�  ���:�  ���;^ :���R��z� ;  
)���  �� 	�� 	B ���� �� �� ;  ��{H�~ d:^�:�@@Rրz� :� ~����  �� 	�� 	B ��  ���B�!�H�L/�� �� �� ��H�;Lz���> M{7��� I;@  �^@�^HAՀ#�^r| Hbx  � X�� �  ��~��N� AՀ#�b| Hc7  �[ X�w �W  ��~I�N� :� �����- @� �
�{4�:� ��  H  �^
�zz�:� ��  H  � r�� pA݁�8!�� (|��A��N� !        ����#�R�* '�                ��� ������|�� (�!��`\  �A  < D� 3� @| �A݀`}  �|  c~  �| 0;_��;> � r�� (���{5' ꀁx(5 	|�z��b�  c5  �� "c  cC  ~��cb  N�!A݁�8!`� (|���N� !        ����#�R�* )       #�R�* �       T   H �       @    #�R�* 3                �'�p%�c�#���U     (      "  , �  �6    $6    <6    �7    �7    �  � �"    �  � �"    x  t �"    |7    �7    7    �6    6    0     �     �6    �     �     @  < T"    	|     	�6    	�6    	�6    
d6    
�6    �  � �"    �  � �"         #�R�* '        T   H �        �    #�R�* 40                   (        , @       #�R�*         T   H �       p    #�R�* 4�                   ,        0 `  7    T7    �7           ���|�#�j�Va�#�R�* /P       T   H �         �    #�R�* 3�                   0        4      h       D � � � � �  p � � � ( T X ` 	� &� .� /� .� /� . 4<           @  �               L l 9       �      :       
                
                         
                         
                            
                         
                            
         	       
                   h                   �d���aG���%�        �    �                 !     �  U    �                         U    �                         �    �                        �    �                      �  �    �                        U    �                  f      �    �                      �  �    �                      �  �    �                       �                                      �                                                                  ���uE�v1�                }                      ����                                        � �                              �                                   @ �� �                            �                                   @ �� K                                                        ���������a�8���@���H���P���X|�� (�!��`\  �A  < D� 3�  | �A݀`}  �|  c~  �~j- @� ;`  �~hH  $;��cc  c�  K���;`  �~�;` �~�A݁�8!@� (|��a�;N� !    ����#�R�* )�        ��k��� ��.VuA    H  �        @           #�R�* 1    ��                                         C @C 
@C D�C H�C I@C M�C j�C q`C  p                        �  ��                                                                     #�R�*  #�R�* �        #�R�* 8�'7nu "X'7nu $        #�R�* 0P'7nu  �#�R�* 9 #�R�* 9�        #�R�* 3 '7nu  #�R�* +�#�R�* *�                                        -      �   " �    #�R�* 2         ~Ϫ�6 [�                        �������  �uc����.�?�        #�R�* :0#�R�* 5P                                                                                                                                                                                                                                          P                  P    #�R�* �#�R�* 1 #�R�* �#�R�* *X'7nu   '7nu  xC                                     �   9                         8!� �      �    #�R�* /P#�R�* 1 #�R�* /P#�R�* /�                                                  ��c$~�h`O��          @   x                        z��        �    #�R�* ' #�R�* 1 #�R�* ' #�R�* *�                                                          `                           ڲ�/       �    #�R�*  #�R�* 1 #�R�*  #�R�* *�                                                          �  -                         ޯآ  �                         h#�R�* '�                                                                   �                  `#�R�* )�                                          ��8�ѶM,"�LP                                              `#�R�* )                                                                    @                   x#�R�* )�                                                                   `                                         3                  #�R�* �                #�R�* �                        #�R�* �#�R�* �#�R�* p#�R�* �                                        #�R�* 0З_�@ �     7�                                                                        �!�Wp���X�                                                                                        �   �   C r�        C t�        C u�                         000`p00 
 %��������@@@@@@@@@@@@@@@@@@@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@                  0                             �                       @       (     x       @     �       `     �           �            �      8     $   �                                0              H              X              h         ��?=�L��:                   (             @          P                l            4             l                                                                                                                                                                                                                                                                                                                                                                                                                     ��s��lo
߂�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��s�Xo   6�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   7   " �  #�R�*        '7nu                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ��qҳ����Y7 (                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��s�Xo   7@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   7`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   7�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   7�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   7�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   7�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ��s�Xo   8    p            #�R�* �#�R�* �        #�R�* #�R�* �        #�R�* |#�R�* � BA    #�R�* �#�R�* 8#�R�* � BA    ��������@@����������\����@@@\����@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�����������������������������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����������������������@@@@�������@@@��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ¥"�:��ܛ?�e@@@@@@@@#�R�* 4#�R�* � BA    #�R�* &�#�R�* �       #�R�* &�#�R�* � BB                                                                                                                                                                                                                                                                                                                                                                                                                                                     ��ƃ;���hC�}�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ĉs�Xo   8�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ŉs�Xo   8�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   Ɖs�Xo   8�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ǉs�Xo   8�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ȉs�Xo   9     t                                                             �        
                                          <          	       B1                      B2              �               ������   	\����m���   \�����m�������   ��������   m����m����m�   m����m������m����   
m����m����   m����m������   m����m�m������m�   m����m�m��m�   m����m�m�����m�   m����m���m�����   m����m����m��m�   m����m����m��m�   m����m����m�   m����m���m���m�   m����m����m���   m����m���m�����  ɦn"k0���Z������   �@��@��ą�����ň   �@��@���È   �@��@������������ɕ��   �@��@���ŗ����            '7nu "�'7nu #�                                                '7nu #�                              U                     �        E   !         U   �        j   �         �         "   �         $   �         %   �   �     '   �         )   �         0   �         2           �  C         �  W         �  g   �     �  �   �                       9                ʇ���5��{��i           
           '7nu $�'7nu %         '7nu %�                        '7nu %                         ;��:���  �  (                           h             �                                                                                                               �                p   �   `                                     �             @  `               	�  �  	@             �     `           �                P  	          `  
0         p  �      �^n�^`�n��d     �  P         �  p         �  �         	P            	`   p                                                                                                                                                                                                                                                                                                                                                                                                                                                      ̉���^�_�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ͉s�Xo   9�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   Ήs�Xo   9�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ωs�Xo   9�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   Љs�Xo   :    @�  #�R�*                   D                  	       B1                      B2              �      c                      D                E                F                G                H                I                O                                P             !   Q             "   R             #   T             $                %   X             &   \             '   `             (   d             *  p             +  	   ��WQ(��b_�             ,  
0             -  �             .  P             /                0  �             1               2  0             3  @             4  P             5  `             6   l             7   p             8   t             9   x             :   |             ;   �             <  p             =  �             >  �             ?  0             @  P             A  p             B   �             C   �             D   �            ғ%R�`I,.c�k   E   �             F   �             G  �             H  �             I  �             J  �             K  �             L  �             M  �             N                O  �             P   �             Q   �             R   �             S   �             T   �             U   �             V   �             W                �  m             �               �                 �               �                �                    Ӌ-P.���P�L�           0                             @                          	  0               �               �               �              P              �              P              P               �                                            `              p            *                +   @          ,             -              .   0          3             4   0            5  �            6  ԓx��`�9���v   @            7  �            �                            ��������@@@@@@@@@@@@@@@@@@@@@@�        �                                                               �                                                   I ��                           %00         
                                                                                                                                                                                                                                       ՘B������/��                                                                  :4     �����                                           V  �            0           F                                                                                                                                                                                                                                                                                                                                                   �Iq�fV��i�]�                                                                            	 H                        	 H                                                                                                                                	                   p � �                                                                                     p � �                     p � �                     p � �                     p � �                     p � �             ׉f�<dޤ`�>P          p � �                     p � �  	                   p � �                     p � �                     p � �                     p � �                     p � �  	                   p � �                     p � �                     p � �                     p � �                     p � �                                             �        x � �                     � � �                      � � �             ؈����V��Ck�C   �        � � �             0        � � �              �        � � �              @        � � �                    p �                        � �                      � �  	                   p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p � �  	                   p � �  	           �G� ��F&��          p � �  	                   p � �                      p � �                      p � �                      p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p � �             ڀ�f�w��`�C�          p � �                     p � �              H       p � �                     p � �                     p � �              
       p � �                     p � �                     p � �              
       p � �                     p � �              �       x � �                                                                                                                                                                                ۀ^���zͪo                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ܉s�Xo   ;�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ݉s�Xo   ;�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   މs�Xo   ;�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ߉s�Xo   ;�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   <                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo   <                                                                                                                                                                                                                           W   m          x @ �                                                                                                                                                                                                                                                                                 �Y|� @<A                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �s�Xo   <`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   <�                                                                                                                                                                                                                                                                                                                                                                                          W      c       x @ �                                                                                                              ��_��3���           � �  	                  � � �  	                   � � �                                              F       p � �                         	              F       `   �  	                    x � �  	                   p � �                     p � �                     ` � �                     ` � �                     ` � �                                              
       ` � �                 
    h � �             ����]�X�Xxr�          h � �              �       ` � �              �       ` � �                     ` � �                           0                         0                    � � �              
       ` � �                      ` � �                      ` � �    �         /     �                                                                                  ` � �                       ` � �                             U        ��k�%�JO��   /                                        U          /                                           �      "   /                                          �      $   /     �                                                              �      '   /                                          U      )   / f                                                       	    p � �  	                  p �                      p �              肥1pB�B»��t          p �                      p �     �      0   /     �                                     �      2   /     �                                    	                  @ � �                     p � �                     p � �                     p � �                     p � �                           H                        	 H                                                                                                   �`H(+���                                                                                                                 �                                                                                                                                        �                                                                                                                                                                     �                           �!T,������4                            @                              �                           �                           �                           �                           �                           �                           �                           �                           �                                                                                                                                             d                           �u���;M���-�   e                            f                            y                            z                            {                            �                            �                           �                           �                                                      "�                           '                            �                           �                           �                           V                          �F*�ݒ%�X��64   ^                           f                           n                     ?      v                                                                                                                 
                                                                                                               �                           �                           �                        @                                                   /     ��yՌ3���                              E                           J                           R                           S                           T                                                �     �                        �                                                                                     �                                                                                                                                             ��� �tM"�^���  "�                           a                           f                               F                        @                            E                                                          ��                                                    �                           #)                          �                          �                        @                                                                                    ��F�2�6�aFF  �                                                        c                                                 �                 �    �  �           =� r                       C� r             �                 �    �  �           E� r                       K� r             }            ����      �  �           M� r                       S� r                                        �      �         �    �               U� r                        𘤠^=W�m�vk9  [N #�                        {N #�                                              :    �                     <    �                           �                           #                           �                                                                                                            	                     B    �                      Y    �                           
                                                      �4�h�^Y��  �   
                                                   \                           f                      
    �                          �                      [    �                           �                           F                �      �  �     �    �                         �                                K      �  �                                                                                                            ���ا�����                                                                                                                  P      *                                  3                        W   �   �                        2                           �                        �                                                      	                 *      
      	      	                 
      
                         ������8�     4                       6                       ,                       -                       .                                              5                       7                                              +                     c   2   3   *   +   ,   -   .   0   /   W   �   �                                                    !   "   #   $   %   &   '   (   7   6   ?   @   A   V   4   5  �� HKesDq?�(   Q   8   9   :   ;   <   =   >   B   C   D   E   F   G   H   I   J   K   L   M   N   O   P   1   R   U   T   S     �   �          	    3  *      4  6  ,  -  .    5  7    +   �   p                                    	                                    
     �        �   ����    ������ǉ������@Ö���������@����@`@����������|�����K���������������   	�      �      �      �   ���������������������������������\����@@@\�����@@\����@@@\����@@@\���@@@@\  �϶�T�~�������@@@\����@@@@@@@@@@@��������  ���Ka��������@@    @              @       @      @  @                                                                                                                                                                                                                                                                                             \�@@@@@@@@    ��������@@@@@@@@@@@@@@@@@@@@@@\����@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@                ����������������������@@���������  ���=�h���Τ�\����@@@\����@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�����������������������������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����������������������@@@@�������@@@��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@    ���    ��<    �� @ ��                                                                                   f      j  �  ��j��W���T��   j  �   j  �   g   �   o         o         o         o         j     l����          .        #       =   %   .          >   %   -   Y             =                   �                   �        6     E   %   -   Y         \     6             �        7     E   %   -   Y        >   %   -   Y        5     7             D                        -   H        =        9      ,   `        �   *   3          !   /  �[-�4�{��!�O     �   c                  9        A   %   W   �      !  �   #       4     :         �   #   �      -   [        E        ;     =   %   /   �         \      !  �   #       3     <      !   /   c                  ;      k     l����       j     j     j  !   l����       n BA   o           D   %   -   H        E   #        -   Y        E        =     >   %   -   Y        =   %   -   H        5     =      !   *     �   >   �   *  ��k����#��T}        N   L      N        �   a          
          !   *     �   >   �   *        N   L      N        �   a          
          !   *     �   >   �   *        �   L      N        �   a          
             -   [        E        >     >   %   -   [         	     ?     >             =         
     ?         	        O   %   *            
        P   %   *           =   #   6     A   %   W            W   m        F         i  ����������t�   "   W   d   q           F   L      N        �   a          
                   i      "   W   d   q           A   L      N        �   a          
             W   �        F         j     X   %   /   �               j        A   %   W   �              E               W   m        F              E   #               X         /   �        �   
     @      /   �        �        A      /   �          2   �        M        B     �E��x�Ȧe^�   /   �          2   �      !  �   *   2             /   �          2   �           B         5        A        @         /   �      #   7   j  #   l����          /   �          2   �      %   .   p         /   �          2   �        M        C      /   �          2   �      !  �   *   2            C      c                  k  #   l����          5         Y         /   �      #   7   !   /     M   c  %                               R   %   *     �7���Q�61�H                  W   m        F              S   %   *                          T   %   *         n      l����       o         !       �   L      L        =      ,   `         K      *   3            >   %   -   p        �   %            !          %   -   \   	   "   -   f   �   -        N   L      N        �   a          
                j  &   l����       j  (         c                     k  (   k  &   l����          ,   `     �F6���!\x�ә       �            C        D     D   #   7     E     D        =   #   7     E              �            o                 F   n      l����       o            �     {               *              D   >   q           �     �   a         
                o               n      l����         G     F      n      l����         =   #  *   n      l����       o         !       �   #  ,   #  +           H        ,     �   
     ���;�e�Ӊ�3�  I     +     ,   >       3            �        I     ,     �   /   #  ,     H     I              +   q            �   q                  #  +              �     ,        J     �   #  .     K     J        ,   #  .     K              .   #  -     -   L      a                     +     -   >   q           �     -   4   L        �      a         
          p  ,         o                 G      n      l����         �(w�M9�h�V  =   #  *   n      l����       o           �   #   �         o               l����          	              Q   %   *         l����                Z      c                     5               j  /   l����          W   m        F        L           M     L              M                 �   %   /   �                                 /   �        D   	     N     �      /   �           O     �      7        O   !   /     �   c   ���F7�d���m�                  P     O      !   /     �   c                  P        Q     N        =   %   -   H         W   m        F        R     D   %   /   �        E   %   -   [        S     R        =   %   /   �        >   %   -   [        S         /   �         ,   `         K      *   3            Q            k  /   l����       j     l����         3      !     %              �   #   !     �   %   *       
   !   *     �   >   �  xHB$OŊ��~   *        �   L      N        �   a          
            �   #        �   #        �   #        �   #         �   #   "     �   #   7     �   %   -   q        �   %   -   r      !   -     �   >   �   -        �   L      N        �   a          
          !   -     �   >   �   -        �   L      N        �   a          
          !  �   %   .          !  �   %   .   �      !  �   %   .   �        �   %   /   �        �   %   /   �        �  W����y��/W   %   /   �      !   W   q           �   L      N        �   a          
            �   %   W           �   #   (   !     q           �   L      N        �   a          
            �   #        �   #             k     l����       j     l����         4              k     l����       k  !   l����       k     k     o         o                  j  1   l����         E   %   -   [         /   �        �        T      ,   `        �  �BF$>䪟Xl|   *   3            U     T         ,   `        �   *   3            U         [   k  1   l����                n BB      7   #   7      [        5        V     V         e      f     j  �   j  �   j  �   g  3      .          �              =   %   .                       c                    =   %   -   H        E   %   -   [                        e     f      j  �   j  �   j  �   !   /      7   c                           ��~py5v�Li�         e      f      j  �   j  �   j  �   j  �     �   #  �     �   a          �       %  �           �     �   a          �         �   a                 a          �             c  �                        a  8              #  4     @   #  6              6     �              6     4   
         !  5     6   A        M   *  5                         !  5     6   A        6     �   /   a  9                 3          *  5      ?$#��51�t�                 6     �   /   #  6                    5            �   #  7     4   %  7          !  7   c                                 �   a           �       !  �   c  �                 e         h      :                      c       +   P            c                      �                      �       +   0            W       +   @            7       +   �            �       +   �            �       +   `            �       +  q�p��d��E��   �            �       +                �       +   �            �       +   �            �       +   �            �       +   �            �       +   �      
      �       +   �            �       +   �            �       +   �            �       +   �            �       ,   �            �       ,   �            �       ,   �            �       ,   0            �       ,   �            �       ,  
                  ,   �                  ,   �     [�ً�X�H�               ,   �                  ,   �         
         -   H                  -   [                  -   Z                  -   V                  -   0                  -   L         
         .                    .                     .                    .                    /   0            +       /   @            ,       /   P            -       /   `            .       /   �            0       /   p           �J�w�!Y�`�   *       /   �                  /   �                  /   �         
                  �                     �     �                                      
     ;       /               ;       '               E                     I      	               g                
     �              4                             9                 9            E        U        j        x                 �     "   �     $   �     	���������  %   �     '   �     )   �     0   �     2                          -      �     �  C     �  W     �  g     �  �                      ��������@@@@@@@@@@@@@@@@@@@@@@�                                                                                                                            |   ��                                                                       ��0                                                                                                      
���k(��k�                                                                                                                                                                  P                                                                       
                                             	                        	               
                                                                  
               :                  $             �v��|�E��@     X  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �s�_��  W
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   A�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   A�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   A�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   B    � #�R�*         ���V  )^ʷ�        �쯉�                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ��5�O�h�ݔ                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �s�Xo   B@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   B`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   B�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   B�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   B�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   B�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   C  �����                                  0                                     P  `  P ���������� @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                ��������@@�����@@@@@������@@@@@@@@@@@@@@@            \���@@@@@@@@@@@@@@@@\������@@@@@      �          @@@@@@@@@@@@@@@@@@@@@�@@@@@@@@���������������������������������������������������@@@@��������@@�������@@@@@@@@@@@@@@@@@@                                @@                      �       �          ������@@@@����@@@@@@          ������@@@@@@@@@@  �l==�w/i;��������@@@@����@@@@@@           D�����9{���.���������@@����@@@@@@   ;       ��������@@@@@@@@                                                                                                                                                                                                                                                                                                                                                                                                                                  _�����D��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �s�Xo   C`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   C�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   C�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   C�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   C�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo   D    8� #�R�*         쯉�  �   `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           !�BE�n]��ZT @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "�s�Xo   D@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   #�s�Xo   D`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   $�s�Xo   D�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   %�s�Xo   D�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   &�s�Xo   D�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   '�s�Xo   D�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   (�s�Xo   E                                  ���@⨔���@あ��       �  E�   @  2  
�   T  �  `            ���� � �� \���m�� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \�  )�͐b��vk+���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���  *u
F{��m5L�� \���� \���� \���� \���� \���� \���� \���� \���� \���� ��������@@                     �������� \�� m����m����m���� m����m������m���� ������ ����                                         �                       ����                  �                      ����                                        ����                  @                       ����                  p   @                                        �                    
                        �                                   +��
����&�                                  	                  0                        
                  `   0                                      �   @                                      �                                            �   �  �                                                                                P                                           �                                            �   @                	                        �                     ,��Qw%j&KA��	                                           	                        @                    	                        p   @                                        �                                            �   @                
   ����                  	                                            	0   �   �      �                           	`  0  0      �                            	�     �               ����                  	�                       ����                  	�      -�b�:r>w8P  	�   E           ����                  
                        ����                  
P      	�   G           ����                  
�      
   	�                                
�    
P  �          ����           J          �  �  �  0                           @  @  P  *�      7                     �      D                                       p     �  D   �                           �  �  
�  @   �       ����                         
�   J   W                   .������#�k���                  �  T   �                           0  `  	0  m   �                                   	0  f                                     	`  7               �             �  0  �   �   �            �             �  �  �  �  8            �                0  �  d               �             P  @  �  �  �            �             �    �  �  �            �             �  �  �  �  x            �                     �  �  p      /�w�jB�[m�;�        �                     �  �  �            �                     �  �  �            �             p     �  X              �             �  �  �  
  �            �                     �    �            �                     �    �            �                     �  ^              �             `  p  �  �  �            �             �  �  �  �  P            �             �  P  �  |  @            �             �     0�]��\�m�z�(>  �  p  0            �                     �  j  (            �                     �  v  8            �                     �  �  H            �             �  @  �  �  p            �             �    �  �  `            �                     �  �  X            �                     �  �  h            �                     �  �  x            �             �  �  �  �  �            �             �  `  �  �  �            �     1���]�h�"��&             0  �  �  �            �                     �  �  �            �                     �  �  �            �                     �  �  �            �             �  P  �  �  h            �             �     �  �  �            �                     �  �  �            �                     �  �  �            �             �  �  �  �  (            �                     �  �               �                     �  �  0      2��������6�        �               `  �   R               �             @  �  �  "  �            �             p     �  �  X            �             �  �  �  �  H            �                     �  �  @            �                     �  �  P            �             0  �  �    �            �                 `  �  �  `            �                     �  L               �                     �    �            �             �  @  3�bX��ͪ���  �  �  �            �                �  �  :  �            �             P  �  �  .  �            �                     �  (  �            �                     �  4  �            �             �    �  R              �                     �  @  �            �                     �  �  �            �             p     �    �            �             �  �  �  �  �            �                     �  �  �            �     4�5Ɗ��`��                  �     �            �                 0  �                 �                     �                �             �  �  �   |   @            �             �     �   d                �                 �  �   X               �                     �   ^               �             P  �  �   p   0            �                     �   j   (            �                     �   v   8            �             �  �  �   �   `      5��O��3�*S�
        �               p  �   �   P            �                 @  �   �   H            �                     �  F  �            �                     �   �   X            �             �     �   �   p            �                     �   �   h            �                     �   �   x            �             `  $0  �  �               �             �  `  �                 �             �    �   �   �            �             �  �  6�6�_ҙ�F�9  �   �   �            �                P  �   �   �            �                     �   �   �            �                     �   �   �            �             �  �  �   �   �            �                     �   �   �            �                     �   �   �            �             @  �  �   �   �            �             p  �  �   �   �            �                     �   �   �            �                     �   �   �            �     7���A���U�iv             0  �      �            �                     �   �   �            �                     �     �            �             �  !`  �  l  �            �             �     �  <  @            �             �  �  �  $               �                P  �                �                     �                �                     �                �             �  �  �  0  0            �                     �  *  (      8���_[�S�@���        �                     �  6  8            �              @   �  �  T  `            �              p   �  �  H  P            �                     �  B  H            �                     �  N  X            �             !   !0  �  `  p            �                     �  Z  h            �                     �  f  x            �             !�  "�  �  �  �            �             !�  "P  �  �  �            �             !�  "   9��T�1i���G_E  �  x  �            �                     �  r  �            �                     �  ~  �            �             "�  "�  �  �  �            �                     �  �  �            �                     �  �  �            �             #  #�  �  �  �            �             #@  #p  �  �  �            �                     �  �  �            �                     �  �  �            �             #�  $   �  �  �            �     :��X�Wa�ڈ(                  �  �  �            �                     �  �  �            �             $`  '0  �  ,  �            �             $�  %�  �  �  @            �             $�  %P  �  �               �             $�  %   �  �              �                     �  �              �                     �  �              �             %�  %�  �  �  0            �                     �  �  (            �                     �  �  8      ;���U�l���R        �             &  &�  �    `            �             &@  &p  �    P            �                     �    H            �                     �    X            �             &�  '   �     p            �                     �    h            �                     �  &  x            �             '`  (�  �  \  �            �             '�  (   �  D  �            �             '�  '�  �  8  �            �                     <�Јg��"Y�  �  2  �            �                     �  >  �            �             (P  (�  �  P  �            �                     �  J  �            �                     �  V  �            �             (�  )p  �  t  �            �             )  )@  �  h  �            �                     �  b  �            �                     �  n  �            �             )�  *0  �  �               �             )�  *   �  �  �            �     =��"pHj)z��^�                  �  z  �            �                     �  �  �            �             *`  *�  �  �              �                     �  �              �                     �  �         e                  .  .�  -  /\  3(  3�  2t  4$  4   4H  3�                      0  /�  04  /�  0X      .�  0�  0�  1T  3p  C�                      1  0�  10  0|  1�  1x  1�  4�  4l  C�  -@  .`  .<  .�          2  1�  2,  ,�  7  2�  3  2�  3L                                  4�  >�� l��p�͍  3�  5   4�  5D  4�  5h  Cx          ,h      C�  88  9�  :T  <�  =�  ?d  ?�  B  BX  A�  B�  B�  B�  B|  C0  C  CT                      D  ,|              @              @  ,�              p               J  ,�              �               �  ,�              �              �  -              �              d  -0              �              �  -T                             �  -x              P              �  -�              �              �  -�              �              �  -�          ?��#	�YH�W�      �              �  .                            X  .,              @              
  .P              p                .t              �                .�              �              ^  .�  ,�                         �  .�              0              �  /              `              |  /(              �              p  /L              �              j  /p              �              v  /�                             �  /�              P              �  /�              �  @�U_�>�jV��c;              �  0               �              �  0$              �              �  0H                            �  0l              @              �  0�              p              �  0�              �              �  0�              �              �  0�                             �  1               0              �  1D              `              �  1h              �              �  1�  -�          �              �  1�              �              �  1�  -�                     A�,�P�oZ��uU      �  1�              P              �  2              �              �  2@              �               R  2d              �              "  2�  /                        �  2�              @              �  2�              p              �  2�              �              �  3              �                3<  /8                         �  3`              0              L  3�              `                3�  /�          �              �  3�              �              :  B<��^� �*�[  3�              �              .  4  .�                         (  48  /�          P              4  4\              �              R  4�  -d          �              @  4�  -�          �              �  4�                              4�              @              �  5              p              �  54              �                 5X              �                5|                               5�              0               |  5�              `               d  5�      C���&��a�          �               X  6              �               ^  60  ,�          �               p  6T                              j  6x              P               v  6�  ,�          �               �  6�  6          �               �  6�  2P          �               �  7                            F  7,  2�          @               �  7P  5�          p               �  7t  6d          �               �  7�  5�          �               �  7�  6@                         �  7�              DWi�c:io�]��  0                8  7`          `               �  8(  7�          �               �  8L  7<          �               �  8p  6�          �               �  8�  5�                          �  8�  7�          P               �  8�  7�          �               �  9   6�          �               �  9$  7�          �               �  9H  8�                         �  9l  8�          @               �  9�  6�          p               �  9�  8\          �                 9�  8�          �      E�;�C���j���;           �  9�                               :   8�          0              l  :D              `              <  :h  :          �              $  :�  9�          �                :�  9|          �                :�  8                           :�  9X          P              0  ;  9�          �              *  ;@  94          �              6  ;d  :0          �              T  ;�  :�                         H  ;�  :�           @              B  ;�  9           p              F�5�No�2	�Q�  N  ;�  :�           �              `  <  ;,           �              Z  <<  :x          !               f  <`  ;          !0              �  <�  <L          !`              �  <�  ;�          !�              x  <�  ;�          !�              r  <�              !�              ~  =  ;�          "               �  =8  <(          "P              �  =\  ;t          "�              �  =�  <          "�              �  =�  =           "�              �  =�  <�          #              �  =�  GH�"�0W�a���  ;P          #@              �  >              #p              �  >4  =H          #�              �  >X  <�          #�              �  >|  =$          $               ,  >�  >           $0              �  >�  >h          $`              �  >�  =�          $�              �  ?  =�          $�              �  ?0  <p          $�              �  ?T  =�          %               �  ?x  >D          %P              �  ?�              %�              �  ?�  >�          %�                ?�  ?@      H�^�چ����\      %�                @  ?          &                @,  =l          &@                @P  >�          &p                 @t  ?�          &�                @�  >�          &�              &  @�              '               \  @�  @�          '0              D  A  @<          '`              8  A(  @          '�              2  AL  >�          '�              >  Ap  ?�          '�              P  A�  @�          (               J  A�  ?�          (P              V  A�  @`          (�  I��`){���y���              t  B   A\          (�              h  B$  A8          (�              b  BH              )              n  Bl  A          )@              �  B�  A�          )p              �  B�  A�          )�              z  B�  @�          )�              �  B�  A�          *               �  C   B4          *0              �  CD  @�          *`              �  Ch              *�              T  C�  5�          �              m  C�                             f  C�  -�          0          JP-׫=viZ)e�      7  C�  6�          `               e                                                                                                                                                                                                                                                                                                                                                                                                                                        ���@�� �$                   ����@�����@����@  K�����<t��2Q  H     �               @  �  0  p  �    p����  0\����@@@@@@@@@@@@@@@@@@@@@@@@@\����@@@@@@@@@@@@@@@@@@@@@@@@@\��@@@@@@@����`�@@@@@@@@@@@@@@     %�������������   ����                                            �����@������@@@@      0          @����nnnnnnnn����@����������@      �          �  ����@���@Ӊ�����@剅�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@���a���@@@@@@@@@\�   %@     ������������� լ��������  P  �������������@����@@@     p     H  P����@@@@@@@@@\������@�����@���@����@��������  L��
��r��_9��@�����    \������@@@      \�����@@@@      \��@@@@@@@      ����`��         \������@@@      @@@@@@@@@@@@@�@�@Ć�������M\��]@������M\���]@������M}�����}]@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@@�@�@���������@@M}ǉ������@Ö���������@����@`@����������|�����K��}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@@�@@aa```````````````````````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@@  M�j���0M."bg�@@aa@ׁ��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@@�@@aa```````````````````````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@@�@�ŕ���ׁ���@@@@@@@��@@@@@@@@@@@@@@@@@@������M}��������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@@�@�@ׁ��@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  N��ֵʺe�@@@@������@@@@@������@@ @@@@@@@@�@�ŕ���ׁ���@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@@�@�@ׁ��@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@\@���@����@����@��@�������@�������@���������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@ć�����@@@@@@@@@@@��@@@@@@@@@@@@@@\@@@�������M}������}]@@@@@@@@@@@@@@@  O����?�[u)�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@���ĉ�@@@@@@@@@@@@@@@@@@@@@@@@@@\@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@���≩�@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@���ĉ�@@@@@@@@@@�@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  P��c��BN�?T@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@@@@@@@@@aa@���������@���@�������@���������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@@��@M������Ml����Mä����]z@l����M������]]@~@\����]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@@��@@@ׁ��@~@}@}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@@��@@@����  QK��3��)J<�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@@��@@@ׁ��@~@l���Ml����Mä����]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@@��@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@@��@@@\����@~@\��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����  R�j�	W�r�I׸��@@@@@������@@ @@@@@@@��@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@@@\����@���������@����      m����m����m���  m����m����m���  �����@@@@@      @@@@@@          �#:��CK        ������@@@@      \��������@����������@      �        �����  @       �    �  (  �  8  �  H  �  X  �  h  �  	x  
   
�    �     �  0  �  @  �nnnnnnnnnnnn����@����������@      �          ��������@⣁������@剅�@@@@@@  S����_�|M�@@@@@@@@@@@@@@@@@@@@@@@@@@����`�@@@@@@@@@@@@@@\�   %@    	������������� լ��������  �������������@����������@ �   �   	     0����  ��@    BA                                                                      BB   nnnn���@����������@@      @        p  p@@@  �����      nnnn���@����������@@      �   	     �����@@@  @  �                                                      	nnnn���@�����@@@@@@@      X      ��������������  ����  p     �  ThY���Ej�Nk$  p      @������  ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          U�s��n% J��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  V�s�Xo   J�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   W�s�Xo   J�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   X�s�Xo   K    � #�R�*         )^ʷ�  D               �  `                                                                                                                                                                                                                                                                                                                                                                                                                                                                         Y�y!��S�g� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  Z�s�Xo   K@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   [�s�Xo   K`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   \�s�Xo   K�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ]�s�Xo   K�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ^�s�Xo   K�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   _�s�Xo   K�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   `�s�Xo   L                            0     p      0�����@����@�����\���������@@@@@@��������@@�����@@@@@            �������������   ��������        \���         E�                \���     E�  P                                                                                                                  p           7������@@@@\����@@@@@          7����@@@@@@\����@@@@@          7��������@@\����@@@@@                                                                                                            a�ʝ���=��i0�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  b�s�Xo   L@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   c�s�Xo   L`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   d�s�Xo   L�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   e�s�Xo   L�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   f�s�Xo   L�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   g�s�Xo   L�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   h�s�Xo   M  ������������@@@@@@@@@@@@@@@@@@@@@@  �                                �   6 @ @                                                               �a�@������@����������@@@            ���� �s�TU�   �  �     �                                        ��%  �tO �                                                �tO �                                                                                                                                                                                          i��	)0�(IS)�\                                                                                                                                 P  P [�D     @   @ 4��    �  � w���           ��%    �  � :�3
           !N7�           "                                                                                                                                                                                                                                                                                  j�D�\~Ğ��*x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  k�s�Xo   M`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   l�s�Xo   M�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   m�s�Xo   M�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   n�s�Xo   M�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   o�s�Xo   M�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   p�s�Xo   N   ( � [�D   0     ��%  � ��������@@@@@@@@@@@@@@@@@@@@@@�      � @6 �s��ޕ  .�M��           
~6O   [�D       �s����                           �   �                               �                                       �              �ǁ ���        �                                                                                                                       ���� !0                                                                                                        q��R�#��S���                                                                                                                                   /ǉ������@Ö���������@����@`@����������|�����K��                   [�D �       �[�D                                             "                [�D @        [�D  [�D `                [�D �[�D �                                        [�D �                                                   �   X   `   �  �  �  �  �  �  �  �  �  �  �  �  X  r�+��7(d^�  H  h  x  X  �  �  h  �  �  8  �  x  (  H  8  (       �   �                    [�D  ��5���[M��m	H        [�D p������@@@@@@@@@@        [�D �������@@@@@@@@@@        [�D ��������@@@@@@@@        [�D `D�����9{���.�        [�D ���������@@@@@@@@ P@�         ��������@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@ P@�         ������@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@ P@�         ������@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@  s�BU�Р�s�3�@@@@@@@@@@@@@@@@ P@�         ��������@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@ P@�         ������@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@ P@�         ��������@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@�     ,                    	                                  [�D �        [�D p[�D �                                [�D X      �        [�D `  h  @        [�D 	�    �        [�D 
�   �  �        [�D �     P        [�D    t�lm�:�D�  �  �        [�D      �        [�D     0  *�        [�D R     +r                ����@@@@@@      �����@@@@@      �����@@@@@      ������@@@@      �������@@@      m������@@@      mm�����@@@      ��������@@      ���������@      ���������@      ���������@      ���������@      ���������@      ����������      ����������      ����������      ����������      ����������      ����������      ����������      ����������      \�@@@@@@@@                                                    @@@                uD�����K�H                                                                                                                                                                                                                              @@@@@                                                                                                                                     ��������@@��\����@@@@@            @@@@@@@@@@  � ����     @      �                  ���������@�������������  � <� :�   ��  �������@@@@@@@@@@@@@@@@@  v4�)���]�@@@@@@  \����@@@@@@@@@@@@@@@@@@@@@@@@@  ��������@@@@@@@@@@@@@@@@@@@@@@  \����@@@@@@@@@@@@@@@@@@@@@@@@@  ��������@@@@@@@@@@@@@@@@@@@@@@  \����@@@@@@@@@@@@@@@@@@@@@@@@@  ��������@@@@@@@@@@@@@@@@@@@@@@  \����@@@@@@@@@@@@@@@@@@@@@@@@@                                                                                                                                                                                                                                                                                       w��ZUlE�֥w�                        @@                                                        @@@@@@@@@@@@@@@@@@@@            �  �  p  p  �  �  �  �  �  �  �  �  �    �  @  �     �   �  �  )`           (                %m����m���m��������   $                      3                                                                                                                                                                                                                                              x��H)�46�2$�
    �[�D  [�D �[�D �        [�D �[�D 0[�D   [�D 0[�D �[�D "�`  � �                 [�D �[�D �[�D                         �,�K�                                        [�D  [�D"�[�D.@[�DCp[�DB                      �                                                                                                                                                                                                                                                  y�\B�p�y��! `0000    000p`    �� 
 
����                                                                                                                                         �           [�D                                          4��                                          w���                                                                                                                                                                                                                            z`L#�Ⱦ����                                                                                                                                                                                                [�D                                                                                              �                                    �       �       �       �       �       �               �       �       �           4��      �       �       �       �       �       �       �       �       �       �       �     {�pOǗ>d�V	P    �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �   [�D �         ��   [�D �         ŀ     |0����0?:�[�D �             [�D �         �   [�D �             [�D �             [�D �         	    [�D �         
�   [�D �             [�D �         �   [�D �             [�D �             [�D               [�D          #�   [�D          (    [�D          �   [�D          �   [�D          �   [�D              [�D          +    [�D           ,    [�D $         �   [�D (         �   [�D ,  }K�q6T=�`���E         �   [�D 0         �   [�D 4         )�   [�D 8             [�D <         
    [�D @         �   [�D D         :�   [�D H         �   [�D L         �   [�D P         &�   [�D T         (�                                                                                                                                     @ ��                                         K                                      �a��������@@                              ~������ޕ���                                                                                                                                                                                   @@@                                                                       �����������|�� (�!�`\  �A  < T� �!83�@| �AڀSA݁��b (`}  �\  c^  �[
��;
�� �������_���?�����8`  8� K�`w  ����;@  ;  ; ����~��x;@����c�  K��`x  )  A�  �<X:����\Pb�  I�c"  N�!� � P:�  �� `�^ `)� @� ��> P� `~�@A� (�� `z�&�  ��b ~G��rt;>���Ȉ:�  ��  �� H  H�^ `;: {9  �� }9�@@� � �8H  {:$�*�� `z�&�;^�~���Ј� �� �> `;Y {Z  �^ `AՀ#K��h��z��� ����z���! ���z���A ���z���� ���z���� ���&z���^6zw��^Fzr��Vz3��fz0���vy�����y���� x���y���� p���y���� h���y���� `�� ������� P��9��;��;8  ���� �y�' ꀁx(: 	|�z��c  a�  �� ;_������ �{�ꀁ{' ꠁxz�{(9 	|�z�{a�  c  �� "� �� �{�ꠁ{' ���xz��(4 	|�y��c4  c  �� 2���� �{�ꠁ{' � �xz�{(4 	|�{/{a�  c  �� B  �5x��ߝn; k{�� �� �z�����z�' � �xy��(5 	|�{�c.  b�  �� Rꠁ� �{�� �{' ���x{5�(/ 	|�yիb�  c  �� bꀁz��� �z�' ���x{�(5 	|�y��b�  b�  � r���z�����z�' ꀁxy�s(6 	|�z�sa�  b�  � �ꠁzO����zT' ���xzի(4 	|�z��b�  bY  � ����zo����zt' ���xz�s(4 	|�z�sa�  bu  �� ��@�z�� �z' ���x{�(/ 	|�zғbV  b  �� ��`�z.�ꠁz4' � �xz��(4 	|�{3�bn  b/  �� �� ��� xy���@�y�' ���xzX�(7 	|�z��c  a�  �� �� ��� py���`�y�' � �xzy�(/ 	|�z�c6  a�  �� ��@��� hy��ꠁ  ���c��؃3X[y�' � �xz��(4 	|�z2�bX  a�  � ��`��� `y��� �y�' ���xz�(7 	|�zӛbt  a�  ��cC  c�  H�!�!  �Q���<h;��9����`���|�b�  a�  �� 28�  bE  c  ~	�c"  N�!A݁�Aڀc8! � (|�����N� !        ����[�D"         ��� ������|�� (�!�A`\  �A  < D� 3� �| �A݀�b (`}  �\  c^  �^�) A� ;@ �^�;_��cC  c�  H�=H ̋^�)� A� H 	\;@ �^�;@  �^ �_� b� o��B;[ � f{8��8  ��  � �Z ~9�@@� ~8�@:�  A� :���A� :� ���0�?�2-  A� ;@  �_� H  D; ���Fz���Y ��  �� 	�8 }��@@� }��@@�   ��	_�x��!�v;  �� H  :�  ��� �_� .:  A�0;   �> ���z���X cC  K��xy �6 �:� ;   )8 A� }6�@;@ @� ;@  -�  A� D�_� r�� vz���; �� ��� �� �� 
�:  :� �Јb�  :�@@��  H  ���{:��� b�  K��xw �~� �;  ;@  *: A� ~8�@:� @� :�  -6  A� (��Vz���; �� ��� �� �� �:  H  4:�  �� �V{6��[ ��� �� Ē� � �V  ;   �> :�  �� ;   � �_� ��� ����B;[ �� �{7���  �  }��@@�  �7 � �� 
�� 
}��@@� }��@;@  A� ;@��A� ;@ �_�0��2.  A� ;   �?� H  4:� ��F{6��V �  }:�@@� ;  �?� H  :�    �O�A���V�F������ ��� -�  A� @; S�;@J�^;  �>:� ��&:� P�� �;  � ;@ �^$H  �_� ��� ����B;[ �� �{7���  �  �7 �� ~6�@@� ~9�@;@  A� ;@��A� ;@ �_�0��2-  A� :�  ��� H  4:� �7  ���Fz��� }��@@� :� ��� H  :�  ��� �_� .:  A� @; S�>; J�:� ��:� ��&;@ ��^ �;  #�> ;  2�$H  ��Vz���:  � �}9�@@�  �� �� �� �; �}6�@@� }8�@;@ A� ;@  -�  A� @:�J��:�S��;  
�>;  	�&;@ ��^ �:� �� :� ��$H ��V{:���  �� �~7�@@�  � �; ��� �� �~8�@@� ~6�@;@ A� ;@  -:  A� @; J�>  ��,"֕Z棉��; S�:� ��:� 	��&;@ Ƴ^ �;  �> ;  
�$H ��_�� �� ���B;[ ��� �z���  ��  �� �� }��@@� � �� }��@@� }��@;   A� ; ��A� ;  �?�0�_�2.  A� :�  ��� H  D:� ��F{6��V ��  � �7 }:�@@� }8�@@� :� ��� H  :�  ��� �� -�  A�L�F{:���  �� z�C,b�  � �Hj� 9�| Hb�  K�`z  V4Ј���6{7���  �W z�C,cV  � �HkY 9�| Hb�  K�`w  ~�4�����&{:���  z� b�  ꠁHj� �| Hb�  K�`y  :4Ȉ�^�z����  z� b�  � �Hj� Z�| Hb�  K�`t  ~�4����&�{:���  ��   �7~%��L�>�z�C,b�  ꠁHj� �| H~� �;@ N   A� ~:�@:� A� :�  -6  A� D��z���� b�  K��xy �{: ȈcC  K�`v  ~�4���� �H  L:�  �� ��z���8  �X {:C,cT  ꠁHkV ~֨| Hb�  K�`w  ~�4��� �;   �> ��z���V  cW  � �HkY 9�| Hb�  K�`t  ~�4���� ��{6��V  cW  ꀁHkU ~��| Hb�  K�`x  4���>$:�  �� ��z����  � ��: �� �}��@@� }��@:� A� :�  .4  A� ��6z���  �� {C,b�  � �Hj� ~��| Hb�  K�`u  ~�4���^�F{4���  �� z�C,b�  �@�Hj� �| Hb�  K�`y  44Ȉ��  ��2��㡉��W:�  �� ;@  �^ H  �;�P:� T���b�  ;   �6  �6 :� d���b�  ;@  �T  �T :� y���b�  :�  ��  :�@�@�z�' � �x(4 	|�{�cX  b�  ��r�� ࢻ 貿��:���~ߡ*:� 
����;@  �_�`�_�hAՀ#K���AՀ#K���A݁�8!�� (|���N� !        ����[�D�x                        �����������|�� (�!��`[  �A  < D� c�  ;��?� ��A݀�B (`|  �;  c>  �>�) A�  ;  �>�;=P?9 c#  cb  H�H ؋>�)� A� H �;  �>�;   �> ;<  ���?  ����{6����{5' ꀁxz׻(5 	|�z��b�  c5  �� r:� d��  �=  *9  @� �>� ~��� v{4���    �BSѢg����L�) @@� h>� �� vz��:� �Ȉ���z��ꠁz�' ꀁxz��(9 	|�z��b�  b�  �� r�=  :� ~��| H��  AՀ#K��x�  )�  A� ��  ;  8�| H>� ~��� vz��~�����ꀁz��� �z�' ꠁx{4�(8 	|�z��b�  b�  � ��  *5  @� �>� ~��� �{7���  ) @@� p>� ��� �z��z��:���;9 �Ȉ���z��ꀁz�' ���xz��(9 	|�z��b�  b�  �X ��  ;  ~��| H��  AՀ#K��p>� ~ݪ�V vzx��  �� �=  {7  Ȉ:� b�  c  b�  K�3�]  ~u�Ө��  34 | H�6 ; ��  ��  :V�ꠁzT' � �x(4 	|�{5�b�  bY  � r�� )� e@� >` ~��  �*j6���F��ð:@ e�T  H  >� =�� �  >� ~���w  �}  �]  zT  ��:� ;�c  b�  b�  K�3�=  �W vzv�~��հ�b�  �]  :` e2�| H{6  Ȉ:� @b�  b�  b�  K�#�^�zy�:�  ��  :�  ��0:� ��P�^@�~H�a h�A `� `�! h�7�:��~��*�� `�a h�~$��:^&���bY  :�@@R��z� ��  �� :��Ը�b�  :�@@Rրz� ��  �� ;>P:�P>� ���@�{7' �`�x(7 	|�zr�bV  c7  �� � 8:}P>s �; 0�@�{' ���x(7 	|�zғbV  c  �� ":� �� 0b�  bc  )�b�  N�!`x  c  �A��ʊ�Β�Ϛ����z���3  . @�  ;  � ��� ��� ���ʚ��H  :�  �� �  ��th�� d�PM��� ��z ���ʚ~��A~Y����> �� �-8��:� @� :�  -�  A���� �~�����^�zu�;   �5  ;   �0:� ��P��`�^h�A x�� p>` =�� p� x��:��~��*�A p�� x��$�^:~&���bx  :�@@R��z� ��  �� :���Ȉb�  :@@@RR�zR �W  �W ;P:�P>� ���`�{' ���x(9 	|�zӛbv  c  �� �[ H;=P?9 � @b�  c#  	�bB  N�!`s  bw  �� ��ʊ�Β�Ϛ����{4��T  . @�  :` �~ ��� ��� ���ʚ��H  ;   � ��: ��� ��>ʚ���� -7��:@ A� :@  -�  A�0�^�zv�:�  ��  ;   �0;   �>P�0��8�� ��� �>@ ~}�� ��� ����  �T�f��|�&��; �~��*�! ��� ���$�>:�&���b�  :�@@Rրz� ��  �� :��՘�b�  :�@@R��z� ��  �� ;>P:]P>R �����{4' � �x(4 	|�{�b�  c5  �� :�P>� ;�� �{�ꠁ{' �@�xz��(4 	|�zY�c4  c  �� b�  cb  Hl�:� ~��� �� �:S �Ҙ��� c  ; �Ȉ�� bU  :U Ҩ�B ����ʊ~Β�Ϛ~���z����  . @�  :� �� ��z ��� ��~ʚ��H  :�  �� ��: ��� ��>ʚ��:Z ; �xr� A� �  � ��  �� H  �� �� ;8 ���c3  >� ~��:U �:� �c#  bD  b�  K�3:� ~��:u0Ө��  ��  � 	�� 	B ��;   �> ���z��:�  ��    �b:2�v�p��4�E:`  �~0:� ��P�p�>x�! �� �>� ~��� ��A ��W�:`�~��*� ��! ��>$��;&���c  :@@@RR�zR �X  �X :��ո�b�  ; @@S9�{9 �5  �5 :�P:�P>� ���@�z�' �`�x(8 	|�zr�bX  b�  � � X:}P>s :���[ P� �z�' ���x(8 	|�z��c6  b�  �� "bc  ~I�b�  N�!`x  � ���ʋ>Β�ϛ>����z���S  - @�  :� �� ��� ��: ���ʛ>�H  :�  �� ��� ��z ���ʚ~�� �c  K��xr �~U �:� M�  A� }��@;  A� ;   .9  A����z��;   �  :@  �^0:�  ��P�0�>8�! ��� �>� ~��� ��a ��w�:@��*� ��! ��>$��  ���5�nz���:�&���b�  :`@@Rs�zs �t  �t ;�ظ�c  ; @@S9�{9 �8  �8 :�P:�P>� ���`�z�' �@�x(4 	|�zS�bx  b�  � :�P>� :W�ꠁzS�� �zX' ���x{5�(8 	|�zիb�  bY  � b�  cb  Hh�:` ~i�� �� �:� �ָ�� bS  :S Ҙ�� b�  :� ֨�B ����ʊ�Β�Ϛ����z���3  - @�  ;  � ��� ��� ���ʚ��H  :�  �� ��z ��: ��~ʛ>�:�:] ;  bC  b�  c  K�3:� א�b�  >� ~}�;3 �:� �b�  c$  b�  K�3;  	�:�0Ԙ��  ��  � 	�� 	B ��:�  �� ;   �> >� �:x0ꀁzu' �@�x(5 	|�zT�b�  bw  �� r;:   ��?�q&$28��,��  �Y  }��@:�  A� :���A� :� �� @�� B.  A� >� ~}�;  �3 0H  �:Z >� ~���� vz��;8 ���:` zu��:�  A� 4~���  ��  }4�@@� DB@ � 	�� 	}4�@A
��@� ,:� zxaM   A� 	�~���~�:� }4�@A
��A� >� ~}�;  � 0H  >� ~]�:�  �� 0>� =�� 0-�  A�h?  ~}�:� P��(�Z,��.��  �W �� ;7 ٸ�c5  ; @@S��  � :��Z0��8�� �T  :� 
ՠ�b�  ; @@S9�{9 �5  �5 :� `:@ @�V  ; ذ�c  :�@@��  R���� ��{2�:�  ��  ;   �0;  �>P� �^�A ��� �� ��! ��3�:@��*� ��! ��>$��;&���c  ; @@  ��k��?�Z7gS9�{9 �8  �8 :��՘�b�  ; @@S9�{9 �5  �5 ;P:]P>R ��� �{' � �x(5 	|�z9�c0  c  � :�P>� ;0� �z�' � �x(1 	|�z�c2  b�  �U "� �z�' ���x(0 	|�z�b2  b�  �U 2� �z�' ���x(0 	|�z��c0  b�  � Bꀁ{' �@�x(3 	|�zT�b�  c  �� Rb�  cb  Hn)�>ʊ>Γ>Ϛ>��^�zp��  . @�  :� �� ��� ��� ���ʚ��H  :�  �� ��: ��: ��>ʚ>�:@  �^ �~���
~��|  �~׆|  �~��|  �~�����>"�^�|  �
  {  �����z��:`  �p  :�  ��0:  �>P�^@�H� ��A �>� ~���a �� Ȳ�:��  �L��<-���7�~w�*�! �� ȳ$�>:^&���bV  : @@R�z �  � :w�Ӹ�bu  ; @@S�{ �  � :>P:�P>� ��� �z2' ꠁx(2 	|�z��� � 8:}P>s :W�� 0� �zP' ���x(0 	|�zыb6  bW  �� "�3 0�� 4: 3� 8c$  b�  b  bc  ~��c  N�!`r  bQ  �! ���ʊ�Β�Ϛ����{4��  - @�  :` �~ ��� ��Z ���ʚ^�H  :�  �� ��� �� ���ʛ��! �~9����> �� �-���:  A� :   .0  A�(�^�zu�:�  ��  :�  ��0;   �P�>0�>8�! ��! �>� ~��A Тa زp�:��~P�*� Т� ز�$��;&���c  : @@R1�z1 �8  �8 :��Ԁ�b�  :@@@  �j�?�����#RR�zR �T  �T :�P:�P>� ��ꠁz�' � �x(9 	|�z5�b�  b�  �V ;P? :��� �z�����z�' �`�xz��(5 	|�zy�c6  b�  �� c  cb  Ha	:@ ~I��T �P �:0 �р�� b�  :� Ԩ�� b7  :7 Ѹ�B ����ʊ~Β�Ϛ~����z���  - @�  :� �� ��: �� ��>ʛ�H  :`  �~ ��� ��� ���ʚ��:Z@: �2  �� �� �2 �� �� �0 �0  ; ؀�c  >� ~��:W �:� �c  bD  b�  K�3:� ~��;70ٸ��0  �9  �0 	�9 	B ��:`  �~ >� �:X0ꀁzU' ���x(5 	|�z��b�  bQ  � r;: �r  ��  }��@:�  A� :���A� :� �� @�� B.    �L$T�U]�xY�yOA� >� ~=�:  � 0H  �:Z ?  ~��� vz��; ؘ�:� z���:   A� 4~	��8  �  }9�@@� DB@ �8 	� 	}9�@A
��@� ,:  z�aM   A� ~��8��~���:1 }9�@A
��A� >� ~}�:  � 0H  >� ~ݺ:�  �� 0>@ =��9 0-�  A�h?  ~��: P�z(��,��.�p  �� �� :� ր�b�  ; @@S9��6  �6 :5�P�zX�q �  :� 
׈�b�  :@@@RR�zR �W  �W ;5 `:� @��  :y �Ȉbx  :�@@��  R���� ���z��;   �  :�  ��0:` �~P�� ���� ��� �� �A �U�:���*�a �� ��$�~:�&���b�  ; @@S�{ �  � :��Ԩ�b�  :`@@Rs�zs �t    �����9`����g�t :^P;P? �����zW' �`�x(7 	|�zv�b�  bO  �� :�P>� :�0�`�z' ���x(2 	|�zӛbn  b  �� "� �z5' �@�x(5 	|�zX�c  b3  �T 2���{0' ���x(0 	|�y��b�  c1  � B���z�' � �x(5 	|�{sa�  b�  �T Rb�  cb  HfU��ʋ>Α�ϛ>���z6���  . @�  ;  � ��� ��� ���ʙ��H  :`  �~ ��Z ��� ��^ʚ��9�  �� ;   �> H 8>  ~=�:� :� Tհ�b�  :�  ��  �� 9� dΰ�a�  :@  �N  �N :� y԰�b�  ;   �4  :@� �z' ꠁx(7 	|�z��c  b  �QB��`��h���9��}�y*;  
�1p:�  ��0��8���z' � �x(5 	|�  �Et���06�<Z{�b�  b  �Q�:��9�@@Q΀y� 9� }����  �� 	�� 	B ���� �� �� ;10:�@@R��z� :� ~����  �� 	�� 	B ���� AՀ#K��AՀ#K��A݁�8!`� (|�����N� !    ����[�D۸        ����!���A��|�� (�!�A`[  �A  < D� c�  ;��?� ��A݀�B (`|  �;  c>  �� �>�) A�  ;  �>�;=@?9 c#  cb  Ho]H ��>�)� A� H |;  �>�;   �> �<"
  {8  Ȉ���z��:�  ��  :�  ��0����>��! h�� `>� =��� `�� h���:��~ٹ*�� `�� h��$��:�&���b�  :�@@Rրz� ��  �� :���Ȉb�  ; @@S9�{9 �6  �6 :�
0;<  ���:�    �k�����u/��*8  A� ~���7��~���~���:� @��삞ʊ�Β�Ϛ����z����  - @�  ;  �> ��� ��� ���ʚ��H  :�  �� �� ��� ��ʚ���> �7�Ȉ�"~������{6�:�  ��  ;   �0;  �>P�P��X�� x�� p?  =��� p�� x���; �~��*� p�� x��$��;&���c  :�@@R��z� ��  �� :���Ȉb�  ; @@S�{ �  � ;>P:�@>� ��� �{6' �`�x(6 	|�zx�� �� h:}@>s ;<  ���� `ꀁ{2��@�{1' � �xzT�(1 	|�z�b�  c1  � 2b�  b�  bc  	�b�  N�!`r  bY  �! ���ʊ>Β�Ϛ>����z����  -� @�  :` �~ �� ��Z ��ʚ^�  �0a�����A�H  :�  �� ��: ��� ��>ʚ���! �7�Ȉ>  ~���� ��|"� �~8� :@ @� :@  -2  A�$��z4�:�  ��  ;   �>0:�  ��P�0�~8�a ��� �?  ~]�� ��! ��2�:��~�*� ��! ��>$��:�&���b�  :�@@R��z� ��  �� ;�ؐ�c  : @@R�z �  � :�P;=@?9 ��ꀁz�' ꠁx(3 	|�z��b�  b�  � :�@>� ;��`�{����{' � �xzӛ(4 	|�z3�bt  c  �� b�  cb  HV):  ~	�� � � c  ; �Ȉ�� bV  :V Ұ�B ���~ʊ�Β~Ϛ����z6��6  -� @�  :� �� ��� ��z ���ʚ~�H  :�  �� �� ��: ��ʚ>�:�p��x  ���e�T7��g&�s2 A� �  � �  �� H  �V �] :� ��b�  >  ~=�;  �b�  b$  c%  K�3;  	�c�  :� �ֈ��u  �v  �u 	�v 	B ��:@  �^ ��,
  >  ~���4 ��|  �
  {  ���>,:�  �� H >` ~��:U: TА�b  :�  ��  �� ;2 dِ�c8  :   �9  �9 :� y֐�b�  :�  ��  :�@� �z�' � �x(8 	|�z0�b  b�  �2�Z��z��u�:�~~U�*:� 
��`:   �5 �5(� �z�' � �x(9 	|�{�b  b�  �U�:�  �� �:� �: @@R1�z1 ;  )��6  �6 	�6 	B ���6 AՀ#K��|AՀ#K���A݁�8!�� (|����N� !        ����[�Dވ                          �����J�:T�����������|�� (�!�a`[  �A  < D� c�  ?� ;�� ��A݀�B (`|  �;  c>  �>�) A�  ;  �>�?= ;9��c#  cb  HhH Np�>�)� A� H O�;  �>�;   �> ?  =�; ��������� ��  :� 	���b�  ; @@S�{ :� >~���  � 	� 	B ��� � � � :� ?~���� ����; ��Ȉ:���Ȉ� c  ; ذ��� b�  :� ט�B ���^�zv�:�  ��  :�  ��0:@ �^P�~���� h�a `�� `�� h���:@�~ّ*� `�a h�~$��:�&���b�  :@@@RR�zR �T  �T :y��Ȉbu  :�@@Rրz� ��  �� :^P>� :�����ꠁzV' �`�x(6 	|�zu�b�  bQ  �   ��l�pD,M��>� :օ�:` ?~i����� ":Y��Ȉ:6  Ѱ�� bP  :P Ҁ��� b3  :3 ј�B ��8� 	b�  cb  K��Y�>ʊ~Γ>Ϛ~���z����  . @�  ;  �> ��z ��� ��~ʚ��H  :�  �� �� ��� ��ʚ��>� �:8 ��Z��:��Q  �1 :q ӈ�bt  :�@@R��z� :  ?~	���  �� 	�� 	B ���� :� ?~���� ���	�:X ����;8	����� bT  :T Ҡ�� c5  ;5 ٨�B �����z��:�  ��  :�  ��0:  �>P������ x� p�� p�� x���:`�~��*� p�! x�>$��:�&���b�  :�@@R��z� ��  �� :�����b�  : @@R1�z1 �7  �7 :�P> :����ꠁz�' �`�x(6 	|�  ������&~h;E�zu�b�  b�  �� >= :1��:` ?~i��	��� ":�	����:�  ֈ�� b�  :� ׀��� b�  :� ֘�B ��8� b#  cb  K��I�ʊ~ΓϚ~���z���0  - @�  ;  � ��z ��� ��~ʚ��H  :�  �� �� ��: ��ʚ>΃>,
  2�Ȉ:�ВV  >� �:x �>��@b��@z��f���b��%��  :� ՘�b�  : @@R1�z1 ;  ?)��5  �5 	�5 	B ��:@ ?~I��� ����:� ����:x����� b�  :� �Ȉ� bu  :u Ө�B �����z��:�  ��  ;   �>0:  �>P������ �� ��� ��� ����:@�~��*�! ��! ��>$�>:�&���b�  :�@@R��z� ��  �� :�����b�  : @@R1�z1   �� ��Gxl�)�7  �7 ;>P> :����ꠁ{6' �@�x(6 	|�zU�b�  c7  �� >= :1��:@ ?~I������ ";8����:�  Ո��� c0  ;0 ـ��� b�  :� Ր�B ��8� b#  cb  K���ʊ^ΓϚ^����z���0  -� @�  ;  � ��Z ��� ��^ʚ��H  :�  �� �� ��: ��ʚ>�>` ~��:� ��: �� ��5  � :U Ҩ�bV  :�@@R��z� :  ?~	���  �� 	�� 	B ���� �� :  ?~)��T ��T�;4 �٠�;�ؠ��� c5  ;5 ٨��� c  ; ؀�B ����z3�:@  �S  :�  ��0:� ��P����� ��� ��! ��A ��T�:`�~4�*� ��� ���$��:&���b  :@@@RR�zR �P  �P :4�  ��7}�b �sV�Ѡ�b3  :�@@R��z� ��  �� :�P>� :օ����@�z�' �`�x(0 	|�zr�bP  b�  � >� :���:` ?~i���� ":��ՠ�:W  Ҹ�� b�  :� հ�� bS  :S Ҙ�B ��8� b�  cb  K��	��ʊ~Β�Ϛ~���z6���  . @�  :� �� ��z �� ��~ʚ�H  :   �> ��� ��� ���ʚ��� x?= ;9��:Z�� pꀁ|�b�  c�  � "�`�|�bv  bW  �� 2c#  ~��c  N�!ꀁ|�b�  c�  �b:] �`�zW' ���x(7 	|�zӛbx  bY  ��������X��P�:����x�>p:� z����� ��� �>} :s��;>p;P:� ���X� �� �{1' ���x(1 	|�z��b  c/  �� "� �  ��F��o��~��{' � �x(7 	|�z�b.  c  �� 2���z�' � �x(0 	|�z7�b�  b�  �� Bbc  ~��b�  N�!� x>= :1��:�  9���� p�`�z�' ���x(5 	|�zӛbt  b�  �� "���|�b�  a�  �� 2b#  }��b  N�!�`�z�' ���x(/ 	|�zӛbt  b�  ��b:= 0���z0' ���x(0 	|�y�sa�  b7  ����z�����X�~P�����x��p9� y����� ��� ���P>� :����� �ꠁ{3' � �x(3 	|�z�b�  c/  �� "ꀁ{' � �x(3 	|�z�b�  c  �� 2� ��Xz�' �`�x(5 	|�zy�c.  b�  �� Bb�  ~����Pa�  N�!: @�  �  :� Հ�b�  ��  �1 ��  �5 =� ~�z�� @�� H�] L  �!S(��8��"ܑ���W����; :` b  c  be  K�3:0 р�b4  ;7��  �� �� �� �� ��  :P Ҁ�bV  ; �x  �r  :�  Ԁ�b�  9� ���  ��  :� �:  @:�  ; @��b�  �X  �S  �X �S �X �S �X �S �  �  ;5 !٨�c/  9�@@Q΀y� :� =~����  �� 	�� 	B ���� �� �� :  ?~)��W ��W�:� �ָ�;�ظ�� b�  :� ր��� c  ; �x�B ����z.�;   �.  :`  �~0:@ �^P������ ��� �� �� ���: �~��*�! ��� ���$�>:~&���br  :�@@R��z� ��  �� 9��ϸ�a�  :�@@R��z� ��  �� :>P=� 9΅���� �z2' ꠁx(2 	|�z��c2  b3    ��L���q�w���N > :��:� ?~������� ":��ո�:0  р��U b�  :� �Ȉ�Q b4  :4 Ѡ�B ��8� !b  cb  K��U��ʉ�Α�ϙ���^�zw���  - @�  ;  �> �� ��� ��ʙ��H  9�  �� ��Z ��z ��^ʚ~�>� ~��; �:�:   :��Јc  �  �  � � � � � � �  �  � (� (�� 0�� 09� 1���a�  :`@@Rs�zs :� <~���n  �n 	�n 	B ���n �n �n :� ?~��� ���:� �ՠ�9��Ϡ�� b�  :� Ր�� a�  9� ϸ�B ���^�zn�:�  ��  :   �>0:  �P���>��! ��� �� ��A ��T�:`��*�� ��� ���$��:>&���b0  ; @@S9�{9 �1    �� ��7aP"��1 :��נ�b�  ; @@S�{ �  � :~P=� 9΅������zp' � �x(0 	|�{6�b�  bq  � >] :R��;  ?	������ ";4�٠�:r  Ӑ�� c.  ;. �p�� bx  :x ���B ��8� 1bC  cb  K����ʊ�Β�Ϛ����z4��  -� @�  9� �� ��Z ��� ��^ʚ��H  :�  �� �� ��: ��ʚ>�:�  ���?  }��ꠁz��� �z�' �@�x{5�(. 	|�zU�b�  b�  ���:  d� @>  ��x @*3  @� �?  }����z����  ) @@� h>� ~����y��; ؈��`�{�ꀁ{' �@�xz��(5 	|�zS�bv  c  ����� @9� ~/p| H�0 @AՀ#K��p?  ~��� @)�  A� �>@   ���e��X��7��x @:� ~ט| H���y��~�Ј�� �z�ꠁz' �`�xz��(2 	|�zy�c6  b  ���=� }�r�/ @*1  @� �>� ~���U�zp��0  ) @@� p>� ~ݺ���y��{�:���:1 Ԉ��@�z���`�z�' � �xzr�(0 	|�{2�bN  b�  ����� @;  ~8�| H�6 @AՀ#K��h>� ~}���{0�:� �� P:Z�9� @��  ��  �� @:/ �x�2� | H�� Pz�  ��b#  b  b�  K�3� P/��x�� P2T | H�S P9� ��  ��  �� P~/��x�� P2� | H�� P; ���  ��  :S����zV' � �x(6 	|�{.sa�  bW  ���� P� @� @z�  ��bC  a�  c  K�3� @��z9�}٢�Ȉa�  �� @  ��/��a���b:� �}��| Hy�  x�:  @a�  b  c  K�#:3 �ꀁz9' ���x(9 	|�z��b�  b/  ���:� ��� @�� @z�  ��b#  bD  b  K�3� @���z��~���Ȉb�  �� @:� ~.�| Hz0  ��:� @b�  b�  b  K�#:� ?~��� ���9� �Ϙ�:��՘�� a�  9� �p�� b�  :� ՠ�B �����zW' � �x(7 	|�{6�b�  bQ  ��;  �� @� @)�  A� �=� ~�r�7 @:@ ~��| H��z8�~x����ꀁzu����zn' � �xy��(. 	|�{4�b�  bq  ��>@ ~ݒ� @*8  @� �>� }����{.��n  ) @@� p>� ~=����z��z�:���:R Ր�� �z��� �z�' �`�x{8�(. 	|�zx�  �6�.��[ �#��c  b�  ���� @:  ~P�| H�Q @AՀ#K��h=� =z9� ?}���Y��Y!�:���Ȉ;!��Ȉ�� b�  :� ՠ��� c  ; ؀�B ���9 @
  ~/����^�zn�:   �  :�  ��0:� ��P���>��! ��� ��A ��a Ȳy�: �~Y�*�� ��� Ȳ�$��:�&���b�  :�@@Rրz� ��  �� :y��Ȉbr  : @@R�z �  � :�P=� 9΅���� �z�' ���x(6 	|�z�b2  b�  �N > :��:� ?~����!��� ":�!��Ȉ:0  р��T b�  :� �p��Q b7  :7 Ѹ�B ��a�  b  cb  K����ʋ>Β�ϛ>����z���n  -� @�  :@ �^ ��� �� ���ʚ�H  ;   �> ��� ��� ���ʚ��  �������0(�ʅ=� ~}r; ��� Ԋ: ֲ�  �8 :� ���b�  9�@@Q�y� :  ?~	���  �� 	�� 	B ���� �� ;  ?)��� ���%�9� �Θ�:�%�՘�� a�  9� ���� b�  :� Ր�B ����{/�:�  ��  :�  ��0:� ��P�^�>��! ��A �� У س�; �~�*� С� ر�$��:�&���b�  : @@R1�z1 �7  �7 :S�Ҙ�bX  : @@R�z �  � ;>P=� 9����ꀁ{6' � �x(6 	|�z4�b�  c7  �� ? ;��:  ?~	��%�� ":S%�Ҙ�;8  ����� bT  :T Ҡ��� c/  ;/ �x�B ��8� c  cb  K����>ʊΒ>Ϛ����z����  . @�  :� �� �� ��: ��ʚ>�H  :     ���:�	v���rՒ ��� ��� ���ʚ��>` }��:� ���P�:T�ZV��  �5 �U :� Ԩ�b�  : @@R1�z1 :  ?~	��4  �4 	�4 	B ���4 :� ?~���� ���)�:o ��x�9�)��x�� br  :r Ӑ�� a�  9� Ψ�B ����z4�:�  ��  :�  ��0:� ��P�^�>��! ��A �� � ��: ��*�� ࢁ 貞$��:�&���b�  ; @@S9�{9 �6  �6 :O��x�bP  ; @@S�{ �  � :>P>� :��������z5' � �x(5 	|�{7�b�  b9  � >� :օ�:  ?~	��)��� ":O)��x�:6  Ѱ�� bW  :W Ҹ�� b0  :0 р�B ��8� b�  cb  K��Ⴞʊ�Β�Ϛ�����z���  - @�  ;  �> �  �R��l��� ��� ��ʚ��H  :�  �� ��� ��� ���ʚ�΁�,
  }��x�9��:n �p��  >  ~]�;2 �? �@c�@{�g��c�%�  :� �Ȉb�  :�@@Rրz� :� ?~����  �� 	�� 	B ��9� ?}��� ��-�9� �ΐ�:r-�Ӑ�� a�  9� Π�� bw  :w Ӹ�B ����z��9�  ��  :   �>0:  �P���>��! ��� �� � ����:���*�� �� ���$��:>&���b0  ; @@S9�{9 �1  �1 :��א�b�  ; @@S�{ �  � :�P>� :օ������z�' � �x(0 	|�{/{a�  b�  � >� :���;  ?	���-��� ";2-�ِ�:�  ՠ�� c/  ;/ �x�� b�  :� ���B ��8� b�    ��W�B���{��cb  K�ڭ��ʊ�Β�Ϛ����z2��  -� @�  9� �� ��� ��� ���ʚ��H  :�  �� �� ��: ��ʚ>�>@ �:x ��� ��� ���  �� ;3 ٘�c/  :�@@R��z� :� ?~����  �� 	�� 	B ���� �� :� ?~��� ��1�:X ����9�1����� bS  :S Ҙ��� a�  9� �x�B �����z��:   �9  :   �09� ��P�~�����a � �����:��~��*�! �!�>$�>:&���b  :�@@R��z� ��  �� :x����bv  :�@@R��z� ��  �� :�P?= ;9����� �z�' ꠁx(/ 	|�z��b4  b�  �� > :��:� ?~����1��� ":x1����9�  π�� bq  :q ӈ��� a�    �s��jR�-�]9� �ȈB ��8� b  cb  K�ؙ��ʊ�Β�Ϛ����{1���  . @�  :� �� �� ��� ��ʚ��H  :�  �� �� ��: ��ʛ>�>  ~��9� ��ZX��`�zd��f�� �n �� �N  : �p�b  :�@@Rրz� ;  >	���  �� 	�� 	B ���� �� ;  ?)�� ��5�9� �Ϩ�:u5�Ө��� a�  9� Ϡ��� br  :r Ӑ�B ����{.�:   �.  :   �0:@ �^P�������������; �~��*�!����$�>:&���b  :�@@R��z� ��  �� :��Ԩ�b�  :�@@Rրz� ��  �� ;>P=� 9΅���� �{2' ���x(2 	|�z�b6  c7  �� > :��;  ?	��5�� ":�5�  ���9:�n3]3N6Ԩ�:P  Ҁ��� b�  :� Ԉ��� bN  :N �p�B ��8� b  cb  K��u�>ʋΓ>ϛ���z5���  - @�  :� �� ��� ��: ���ʛ>�H  ;   � �� ��: ��ʚ>�>� }ݪ:n ���h�Zp��t�S �� ��  :� ט�b�  ; @@S9�{9 ;  >	��7  �7 	�7 	B ���7 �7 �7 :  ?~	�� ��9�:� ��p�:N9��p�� b�  :� ՠ�� bO  :O �x�B �����z��:   �3  :   �09� ��P��>��!(�� � ��(���:���*�! �a(�~$�>:&���b  ; @@S9�{9 �0  �0 :���p�b�  ; @@S�{ �  � :�P>} :s����� �z�' � �x(/ 	|�{1�b8  b�    �P�K��>�|�S� > :��:� ?~����9��� ":�9��p�9�  π�� b�  :� Ԉ�� a�  9� Ϙ�B ��8� b  cb  K��U��ʊ�Β�Ϛ����z.��n  -� @�  ;  �> �� ��� ��ʚ��H  :�  �� �� ��: ��ʚ>�=� ~}r:S ��� ԉ� ֲ�  �� :� Ԑ�b�  ; @@S�{ :� ?~���  � 	� 	B ��� � :� ?~��� ��=�9� �Θ�:�=�՘�� a�  9� �x�� b�  :� Ր�B �����z��:   �4  :   �0:@ �^P���>��!8��0�0��8���:���*�!0��8��$�>:&���b  ; @@S9�{9 �0  �0 9��Ϙ�a�  ; @@S�{ �  � :�P>� :������ �z�' � �x  �GL �/E't��(2 	|�{1�b8  b�  � > :��:� ?~����=��� "9�=�Ϙ�:P  Ҁ�� a�  9� ψ�� bT  :T Ҡ�B ��8� b  cb  K��A��ʊ�Β�Ϛ����z3���  . @�  ;  �> �� ��� ��ʚ��H  :�  �� �� ��: ��ʚ>�>` ~��:� ���P�ZT��V��  �U �� ;5 ٨�c8  :�@@R��z� :� ?~����  �� 	�� 	B ���� :  ?~	�� ��A�:t �Ӡ�9�A�Π��� br  :r Ӑ��� a�  9� �x�B ����{5�:   �5  :   �09� ��P�^�����H�A@��@�H��; �~��*�!@��H��$�>:&���b  :�@@R��z� ��  �� :T�Ҡ�bX  :�@@Rրz� ��  �� ;>P  ����"�K���>� :������ �{/' ���x(/ 	|�z�b6  c7  �� > :��;  ?	��A�� ":TA�Ҡ�9�  π��� bQ  :Q ҈��� a�  9� Ϩ�B ��8� b  cb  K��)�>ʋΓ>ϛ���z����  - @�  :� �� �� ��: ��ʛ>�H  ;   � ��� ��� ���ʚ�΂>,
  ~7���9��:n �p���  =� ~]z:� �> �@b�@z�f��b�%�  ;6 ٰ�c8  :�@@R��z� :� ?~����  �� 	�� 	B ��:  ?~)��� ���E�9� �ΐ�:rE�Ӑ�� a�  9� �x��� bp  :p Ӏ�B ����{1�:�  ��  :�  ��0:  �P������X��P�P�X��; �~��*��P�!X�>$��:�&���b�  :�@@  ����E�շ�gbBR��z� ��  �� 9��ϐ�a�  :�@@R��z� ��  �� ;>P>= :1�������{0' ꠁx(0 	|�z��b�  c5  �� >� :օ�;  ?	��E�� "9�E�ϐ�:  а�� a�  9� ϸ��� b  : Ј�B ��8� b�  cb  K����>ʋΓ>ϛ����z���2  -� @�  :� �� ��� ��: ���ʛ>�H  ;   � ��� ��� ���ʚ��>@ ~=�:q ��� �� ���  � 9� Ϙ�a�  :�@@R��z� ;  ?)���  �� 	�� 	B ���� �� ;  ?	��� ���I�:Q �҈�9�I�Έ�� bP  :P Ҁ��� a�  9� Θ�B ����{/�:�  ��  :�  ��0:` �~P�����h�`�`�h��; �~��*��`��h��$  ���)�g�r��~��:�&���b�  :�@@R��z� ��  �� :�Ј�b  :�@@R��z� ��  �� ;>P=� 9�������{3' ꠁx(3 	|�z��b�  c5  �� >� :օ�;  ?	��I�� ":I�Ј�:v  Ӱ�� b  : и��� bo  :o �x�B ��8� b�  cb  K���>ʋΓ>ϛ����z����  . @�  :� �� ��� ��: ���ʛ>�H  ;   � ��� ��� ���ʚ��>  }��9� ��Zx�z��n �N  : �p�b  :�@@R��z� ;  >)���  �� 	�� 	B ���� �� ;  ?	��� ���M�:/ ��x�:oM��x�� b2  :2 ѐ��� bn  :n �p�B ����{0�:�  ��  :�  ��09� ��P�^����x�Ap�p�x��  �u����1��S�h; �~��*��p�x�$��:�&���b�  :�@@R��z� ��  �� :O��x�bX  :�@@R��z� ��  �� ;>P> :�������{.' ꠁx(. 	|�z��b�  c5  �� >� :օ�;  ?	��M�� ":OM��x�9�  ΰ�� bW  :W Ҹ��� a�  9� ΀�B ��8� b�  cb  K��̓>ʋΓ>ϛ����z���  - @�  :� �� ��� ��: ���ʛ>�H  ;   � ��� ��� ���ʚ��=� ~z:p ��:������ �3  :S Ҙ�bU  :�@@R��z� ;  >)���  �� 	�� 	B ���� ;  ?	��� ���Q�9� �π�9�Q�΀��O a�  9� ψ��N a�  9� Ψ�B ����{4�:�  ��  :�  ��0:� ��P�>�~��a�  �����{3 �!��A�����; �~P�*��������$��:�&���b�  :`@@Rs�zs �v  �v :0�р�b8  :@@@RR�zR �Q  �Q ;>P>� :��������{5' �`�x(5 	|�zw�b�  c3  �T >� :օ�;  ?	��Q��� ":0Q�р�;6  ٰ��Q b7  :7 Ѹ��Y c8  ;8 ���B ��8� b�  cb  K�ǽ��ʊ�Β�Ϛ�����z���  -� @�  :` �~ ��Z ��� ��^ʚ��H  :�  �� ��� ��� ���ʚ��>  �9� �����:��. ��  :. 
�p�b3  :@@@RR�zR :� >~���Q  �Q 	�Q 	B ���Q �Q �Q :� ?~���� ���U�: ����;8U������ b  : И��� c5  ;5 ٨�B �����z��:   �2  :�    �r�AF��-|��0:� ��P�~�������a����������:��}ع*�!��A��^$�>:�&���b�  9�@@Q�y� ��  �� :x����bv  9�@@Q΀y� ��  �� :�P>] :R����� �z�' ���x(5 	|�y�b4  b�  �� >� :օ�9� ?}���XU��V "9�U����:�  װ�� a�  9� ψ��� b�  :� �p�B ��8� 
b�  cb  K�ť�~ʊ^Β~Ϛ^���z����  . @�  :  �> ��� ��z ���ʚ~�H  :@  �^ ��� ��� ���ʚ���o��=� ~r������9� ��A�zq���  ��  }4�@;   A� ; ��A� ;  �0 p� r-�  A� =� ~�r:�  �� `H  l:Z >` ~=����y��� �2  � � ~4�@@� ~0�@  ��QRؗ�I �&g@� �� �� ~6�@@� >` }ݚ:  �. `H  =� =z:�  �� `?  ~�� `-5  A� H:^��������z���  �� �r :2 ѐ�b.  9�@@Q�y� ��  �� �� H  h:�  �� ;>�?  ~�ꠁ{7' ���x(7 	|�zիb�  c3  �P���fy��:� �� @� @{  ��c#  b$  b�  K�3:�  �� :��>` ~]����z�' ꀁx(/ 	|�z�sa�  b�  ��:  � @>  ~���� @)�  @� �>` }����z���.  * @@� h?  ~����z��:2 ѐ��`�z4����z5' ���xy�(5 	|�yӛbx  b9  ���� @:� ~W�| H�P @AՀ#K��p>� }��� @)5  A� �=� ~=r�q @;  �| H���z��~�  ��x���,���B�А�ꀁz�ꠁz' �`�xz��(. 	|�zt�b�  b  ��>� ~���W @)�  @� �=� ~�z�U�zn��  * @@� p>� =���z8�{�:���:� װ����z��ꠁz�' ���xz�{(3 	|�y�{a�  b�  ��� @;  ~ؠ| H�� @AՀ#K��h>@ ~���U�zn�:� �� P9��:= @�  �� � 
�� � 
�  �� @;1 و�2V | H�U Pz�  ��c#  a�  be  K�3�� P}�ψ�� P3 | H� P: ��P  �O  :��� �z�' �`�x(. 	|�zy�c.  b�  ����� P�� @� @z�  ��b�  b$  c  K�3� @�U�zy�}���Ȉa�  �� @:� �~7�| Hz8  ��:@ @a�  bD  c  K�#:u �� �zy' ���x  �v�t�Po�-��Ѓ(9 	|�yЃb  bo  ���:� ��� @�� @z�  ��bc  b�  b%  K�3�U @��{0�}�π�a�  � @:� ~t�| Hzq  ��;  @a�  c  b%  K�#;  ?)��U ��UY�: �Ш�9�Y�Ψ�� b  : и�� a�  9� Π�B �����z�' �`�x(1 	|�zo{a�  b�  ��:@ ��U @� @)4  A� �>� ~=��q @:� }��| H��{2�~�zՐ�ꀁz��� �z�' �`�xz�(7 	|�zt����>� ��8 @)�  @� �=� ~]z���z���  * @@� p>` ~����z4�z��;4��; ������{6��@�{7' ���xzO{(7 	|�y�{a�  c3  �U�� @:  ~��| H�� @AՀ#K��h?  ~��:� ?~���Y��]�  �J�|�`R����>'9�Y�ΰ�9�]�ϰ��N a�  9� ΀��O a�  9� ψ�B ��� @
  ~������{7�:   �7  :   �0:` �~P�^������A����!��6�: ��*������$��:~&���bt  :@@@RR�zR �S  �S ;6�ٰ�c8  : @@R1�z1 �9  �9 :P>� :�����ꀁz' �`�x(2 	|�zt�b�  b  � >= :1��:@ ?~I��V]��Q ":]�а�:�  Ԉ�� b  : и�� b�  :� Ԙ�B ��b�  b#  cb  K��M�^ʊ�Β^Ϛ���^�zw��7  - @�  ;  � ��� ��: ���ʚ>�H  :�  �� ��Z ��z ��^ʚ~�>� =�9� �������У؊�ڳ �� ��  �� � :/ �x�b6    �����V/p�u�f:@@@RR�zR :` =~i��Q  �Q 	�Q 	B ���Q �Q �Q :� ?~��� ���a�; ��Ȉ9�a��Ȉ�X c  ; ؀��N a�  9� �x�B ����z6�:�  ��  :�  ��0:� ��P���~��a�����A��Ȳ�: �~Y�*�����Ȳ�$��:�&���b�  :`@@Rs�zs �u  �u 9���Ȉa�  :@@@RR�zR �O  �O :>P>� :օ������z4' �`�x(4 	|�zw�b�  b5  �� > :��:@ ?~I��Ya��P "9�a��Ȉ:0  р��� a�  9� Ϩ��� b4  :4 Ѡ�B ��8� b  cb  K���~ʊ^Β~Ϛ^���z����  -� @�  :� �� �� ��z ��ʚ~�H  :@  �^ ��� ��� ���ʚ��?  ~��9� �� �  �˫��%�cU��$�: ֳ  �. 9� �p�a�  : @@R�z :` ?~i��  � 	� 	B ��� � :@ ?~I�� ���e�;7 �ٸ�;e�ظ�� c.  ;. �p�� c  ; ذ�B ���^�zo�:�  ��  :�  ��0:� ��P���>��!�����ТAزW�:`�~�*�С�ر�$��:�&���b�  : @@R1�z1 �4  �4 9��θ�a�  : @@R�z �  � :~P=� 9����ꠁzv' � �x(6 	|�z5�b�  bq  � >� :���:@ ?~I��We��T "9�e�θ�:�  ֠�� a�  9� Ψ�� b�  :� �x�B ��8� b�  cb  K��	�~ʊ^Β~Ϛ^���z����  . @�  :  �> �� ��z ��ʚ~�H  :@  �^ ��� ��� ����  �|<��
<�����>� }��; ��:P��T��V�8  �� �� :8 ���b0  :`@@Rs�zs :@ ?~I��q  �q 	�q 	B ���q :� ?~��� ���i�:� ��x�;/i��x��W b�  :� װ��Y c.  ;. �p�B ����z8�:�  ��  :�  ��09� ��P���~��a�����A���: �~O�*���$��:�&���b�  :`@@Rs�zs �t  �t :���x�b�  :@@@RR�zR �V  �V :>P? ;����ꠁz.' �`�x(. 	|�zu�b�  b3  �X >� :���:  ?~	��i�� ":�i��x�9�  Π��V b�  :� ֨��N a�  9� ���B ��8� b�  cb  K���>ʊΒ>Ϛ���z���  - @�  :` �~ ��Z ��: ��^ʚ>�  �s�8�O�R�~I�H  :   � ��� ��� ���ʚ�΁�,
  }��x�;>�:� �Ȉ�  =� ~�r:v �>@�@bR�@zR�fR��bR�%�S  :3 ј�b0  :�@@R��z� :� ?~����  �� 	�� 	B ��9� ?}��� ��m�:� �װ�9�m�ΰ��W b�  :� ׀��N a�  9� Ψ�B ����z4�9�  ��  ;   �>0;  �P��~��a�����A����: �~V�*������$��;>&���c8  :`@@Rs�zs �y  �y :��հ�b�  :@@@RR�zR �U  �U :>P>� :��������z8' �`�x(8 	|�zo{a�  b9  � > :��:@ ?~I��m��� ":vm�Ӱ�:0  р�� bo  :o �x�� b2  :2 ѐ�B ��8� b  cb  K�����ʊ��  ���W��$�x��"��Ϛ����{6��V  -� @�  9� �� �� ��� ��ʚ��H  :�  �� �� ��: ��ʛ>�>� ~]�9� ��� ��: ���  �. :n �p�bo  : @@R�z :� ?~���  � 	� 	B ��� � :� ?~��� ��q�:� �֐�:�q�א�� b�  :� �p�� b�  :� �x�B ����z��;   �3  ;   �09� ��P���>��!�� � �����:��~�*�! �a�~$�>;&���c  : @@R1�z1 �8  �8 9��ΐ�a�  : @@R�z �  � :�P>} :s����� �z�' � �x(/ 	|�z9�c.  b�  �� ? ;��:� ?~���q�� ":�q�Ր�;8  ����� b�  :� ՘��� c4  ;4 ٠�B ��8�   ��)ā�ZH�_o��c  cb  K����>ʊΒ>Ϛ��^�zt���  . @�  9� �� �� ��: ��ʚ>�H  :   � ��Z ��z ��^ʚ~�>� }��:� �����:����� ��  �7 9� θ�a�  : @@R1�z1 :  >~	��.  �. 	�. 	B ��:@ ?~I��O ��Ou�:� ��x�:�u��x�� b�  :� ԰�� b�  :� ո�B ����z.�:`  �n  :@  �^0:� ��P���>��!������: ��*�a����$�~:^&���bW  ; @@S9�{9 �2  �2 :���x�b�  ; @@S�{ �  � :>P=� 9΅����`�z7' � �x(7 	|�{3�bv  b7  �� >] :R��:  ?~	��u�� ":/u��x�:r  Ӑ��� b.  :. �p���   �*p9�V�����~�bp  :p Ӏ�B ��8� bC  cb  K����>ʋΓ>ϛ����y����  - @�  :� �� ��Z ��: ��^ʛ>�H  ;   � ��� ��� ���ʙ��>  ~��:� ����z �:���� ��  �u �5 :U Ҩ�bY  ; @@S�{ 9� =}���  � 	� 	B ��� � � 9� ?}���W ��Wy�: �и�:�y�ָ�� b  : Ј��� b�  :� �ȈB �����y��:`  �x  :@  �^0;  �>P�>����(�! � ��(���9��~�y*�a �(�$�~:^&���bY  :�@@R��z� ��  �� :7�Ѹ�b.  :�@@R��z� ��  �� 9�P? ;�����`�y�' ꠁx(9 	|�z��bt  a�  �� >] :R��9� ?}���y�  ���W}��E��m� ":7y�Ѹ�9�  ϐ�� b3  :3 ј��� a�  9� �p�B ��8� bC  cb  K��m�>ʋΓ>ϛ��^�zw���  -� @�  :� �� ��� ��: ���ʛ>�H  ;   � ��Z ��z ��^ʚ~�>� }ݺ:� �� ԉ� ֲ  �� :6 Ѱ�b5  :�@@R��z� ;  ?)���  �� 	�� 	B ���� �� ;  ?	��N ��N}�:� ��p�:}��p�� b�  :� �x��� b  : а�B ����{1�:`  �q  :@  �^0:� ��P������8��0�0�8��; �~��*�a0�!8�>$�~:^&���bV  :�@@R��z� ��  �� 9���p�a�  :�@@R��z� ��  �� ;>P>= :1�����`�{6' ꠁx(6 	|�z��bt  c5  ��   �����m�4�>] :R��;  ?	��}�� "9�}��p�:�  ֐�� a�  9� Ϙ��� b�  :� ֈ�B ��8� bC  cb  K��Y�>ʋΓ>ϛ��^�zn��.  . @�  :� �� ��� ��: ���ʛ>�H  ;   � ��Z ��z ��^ʚ~�=� ~=r: ���P��T��V��  �� �� :� Հ�b�  ; @@S9�{9 ;  ?	��5  �5 	�5 	B ���5 >@ bR� ~}�9� ?}���� ����9� �ψ�:�И�� a�  9� Ϡ�� b  : Ш�B �����z��9�  ��  :�  ��0:� ��P�>���H�!@��@��H���9��~�q*�A@��H��$�^:�&���b�  ; @@S9�{9 �4  �4 :��׈�b�  9�@@Q΀y� ��  �� :�P>] :R����  ��EЭ���h*� �z�' ꀁx(9 	|�z��c  b�  �� >= :1��9� ?}����� ":��Ԙ�:�  Ո��� b�  :� Ԑ��� b�  :� �p�B ��8� b#  cb  K��5�>ʋΓ>ϛ��^�zn���  - @�  :� �� ��: ��: ��>ʛ>�H  ;   � ��Z ��z ��^ʚ~�9�  �� H X>� ~�9�@:� T�x�b�  :�  ��  �� :/ d�x�b9  ;   �  � :O y�x�bS  9�  ��  :�@ꀁz�' ꠁx(6 	|�z��b�  b�  �b�:�� ���:`�~0�*��(�Z0��2�P�������:��ꀁz�' � �x(9 	|�{���B9� ���:   �0P�0X�`�z�' ���x(2 	|�zӛbx  b�  ��9��:�@@R��z� ��  �� �� :��  �� �4J.Ed��υ9�@@Q�y� :  ~)���  �� 	�� 	B ���� AՀ#K��LAՀ#K��TA݁�8!�� (|�����N� !    ����[�D߸                                �����������|�� (�!�a`\  �A  < D� 3�( | �A݀�b (`}  �\  c^  �^�) A� ;@ �^�;_��cC  c�  H�H & �^�)� A� H ',;@ �^�;@  �^ `   ;^)`� �{X' ���x(8 	|�z��c6  cW  ���;  �+;^ �; @@S9�{9 �:  �: :�  ��|:�8; :;;8�؈;^:�����  ��  �� �� �� �� �� �� ��  � "��  � ":� ǒ�+(�>+?* �A� ���`�d��:�>;@��^ �:������>�- d@� p��0����*�^*��^v:�n  ��'��<���Fb��*; ::��;^:���;������  ��  �� �� �� �� �� �� �:  �� "�8  �� "��|��#H  ����r;@ 
�^��� �:���;>p� ��@�{5' ꀁx(5 	|�z��cT  c5  �� "b�  	�b�  N�!�>��^��^ �>:� I��:�  ���:� �� � �:���;^@�< �ꠁ{T' ���x(4 	|�z��b�  cS  �V "b�  )�c  N�!���� ����-� dA� X�^��^ �� �:��:_� ����< �� �zT' ���x(4 	|�z��c  bQ  � "b�  bc  )�b�  N�!�^ * �:� @� :�  -4  A�!����z��;   �  :   �>0:   �P�~�>�! h�a `� `�A h�_��:�ߺ~��*�� `�� h��$��;&���c  : @@  ��(�%^�(�a�vR1�z1 �8  �8 :� ;0�ـ�c3  ;@@@SZ�{Z �Y  �Y :�P:�� :�#�נ����z�' � �x(2 	|�z6�b�  b�  �W ;��c  c�  H #�`p  b  �A@�>ʊ�Γ>Ϛ����z5���  -� @�  :` �~ ��[ ��� ��^ʚ��H  ;   � ��; ��� ��>ʚ���A@P�Ј�ݐ`   :>)`ꠁz6' �`�x(6 	|�zu�b�  b7  ���:@ �^ ;  �+;> �:�@@R��z� ��  �� ;@  �^|: h:`::;h�؈:�:�����  ��  �� �� �� �� �� �� ��  �Q "��  �U "�+?* �A� �����;���:�>>;@��^ �: ����~�- d@� p��0����>*��*���v:@n~>�*:�:; �:�:���;>�����T    �7�Z��UV�Xp�Y  �T �Y �T �Y �T �Y �  �t "�  �y "��|��#H  @:�  ���:   �>  :@ �^�:���b�  c�  H%��� ��^�-� dA� \���� �� �:��;?� ����� �� �{2' ꠁx(2 	|�z��b4  c5  �� "b�  bc  ~��b  N�!H  |�+C* �A� ;@ �^ H  d:@��^;  �>  :  �>�:���b�  c�  Hy��)�z��:` �t  �)���:  �  ;@ �^�:_��bC  c�  HA�> ) �:� @� :�  -�  A�d:��`:� M��  :v Ӱ�bt  ; @@S9�{9 ;  ?	��3  �3 	�3 	B ���3 �3 �3 :  ?~	���o���;_�`:_��� cW  ;W ڸ��� bV  :V Ұ�B ����{3�:   �3  :   �0:�   ��ř�w��d�_��P������ x�� p� p� x���; ߺ~��*�! p�a x�~$�>:&���b  :�@@R��z� ��  �� :�� ;�ظ�c  ; @@S9�{9 �8  �8 :~P:?� :�#�ֈ�ꠁzp' ���x(0 	|�z��b�  by  � :���:  ?~)������� ":��:t  Ӡ�� b  : Ш�� bq  :q ӈ�B ��8� b�  c�  K�����ʊ�Β�Ϛ����z���1  . @�  ;  � ��� ��� ���ʚ��H  :�  �� ��� ��; ���ʚ>�;?� �@�{:' �`�x(: 	|�zr�bV  c7  ���b:  ��� �� {  ��:�	 c#  b�  b�  K�3�?� �_�fzz�~���Јb�  �� ;  0�| H{5  Ȉ:� @b�  b�  b�  K�#:[��`�(|�bp    �{.g�6︋����bQ  ��r;_ݔ���{X' � �x(8 	|�{6�b�  cU  ���bAՀ#���r| Hb�  �{��2 �  ��~	�N� ��f{:�:� ��  ���fz���T  -2 A�H  \H  X:;��`�(|�bx  b9  ��rAՀ#K��h��o�� ��� �z���P  :@ ~:�|  �~34���p  AՀ#K���;   �?ݖ;  �ݘH  $��ݘ-�  :� A� :�  .4  A� H |��ݔ������b�  �A8�_��_�-: A� �?�-� @� L�| �:��;?� � �ꠁ{4' ���x(4 	|�zիb�  c7  �� "8� db  	�bb  N�!;@ �A8~:�P|  �b4  ��0;  ~��|  �������.7 A� ���-6  @� D� �;��:� �\ ��@�zq' � �x(1 	|�{2��X "8� dc  I�b    �co������ !N�!�0:� ��� :�$-�  z��~7�@� :� Ѱ�b9  �! �ݖ:@ �|  ����_�cP  �(����.5 A� ��-4 @� L�� �:���:?� �\ ��`�z8' �@�x(8 	|�{S�bt  b5  �� "8� db�  ~I�b�  N�!;  �(�P|  �
  �! ;@ ~8�| H�?� �| �:���:�� ~��֠��_� zW  ���� z  ���< �� �{4��@�{0' ꀁxzX�(0 	|�z��� "�@�z��ꀁz�' � �xz��(9 	|�{�bX  b�  � 28� b�  cF  8�  9  b�  ~)�bb  N�!`p  b  ��������-�  @� L�\ �;?��;� �� ��@�{' � �x(5 	|�z:�cT  c  �� "8� dc#  ~��bB  N�!�~�4���ݘ  ���<$"��b*��ݘ.0  :� A� :�  -6  A�\�?ݘ�ݖX�|  �U4Ј��ݖ;   �?���ݖ���@:_� ꀁzS' � �x(3 	|�z�b�  bQ  �݂:� �� �|�c  b�  ���b�_�@-�A� �?�@.9  @� L�� �:��:_� �< �� �zV' � �x(6 	|�{�b  bU  �� "8� dbc  ~)�b�  N�!�_�-: A� �?�-�  @� L�� �;��:_� � �ꠁzT' �`�x(4 	|�zu�b�  bO  �� "8� dc  ~	�b�  N�!�?�@:� W�P|  ��_�@;   �?� ��@
  z�  ��:_�0�݆z��bC  a�  be  K�3���@
  �� ~p| H�� ~�r֐�b�  ��fz:��:  �6  �� 2� | H��� 9� ϸ��`�y�����y�' � �xyӛ(2 	|�z�  �صU�0���rPbp  a�  ��b�_�@
  �?�
  ~��| H
  ���@��@.4 A� d��@:� �P|  �
  ���fy��bS  {  ����@
  �݆z��:��ЈbC  c$  b%  K�3��� ~��| H��� ��� ��� 9�� �`�y�' ꠁx(4 	|�z��bx  a�  ��b�� )0 @� ;@ �_�PH  �_� �_�P�?�P�?� ��� z�  ��9��0:�� b�  a�  b�  K�3�� ���fy��3�٘�c8  �� ;@ ~P�| HzQ  ��:� @c#  b�  b%  K�#��ݖ:� }Ծ|  �}�4p���ݖ:�  �� AՀ#K��l:`  �~ AՀ#K���;� �@�{' �@�x(0 	|�zZ�cP  c  ��b;  �?� ��� )�  A� ���� :� }Ը| H��fz��~or�x��@�zx��@�zq'   �Z�;p��z�h� �x{R�(1 	|�z��_݂�?� *9  @� t��݆z����  ) @@� `��݆y��{�:8��;Z �Ј� �z3��@�z9' ���xzP�(9 	|�zЃ�݂��� :� ~��| H��� AՀ#K������fy��;_�`�`�{R' � �x(2 	|�{3�bp  cQ  ��b��� ��� ��� z�  ��cC  c  b�  K�3�� ���fy��2�ِ�c3  �?� :  ~р| Hz�  ��;@ @c#  cD  b�  K�#;  ?	����o����:��`:����T b�  :� Ԁ��U b�  :� Ո�B ��:�� � �z�' ���x(: 	|�z��c.  b�  ���b;  �� �?� )�  A� ��� :` ~S�| H���fz��:��Ј���{.�� �{1' ꠁx{{(1 	|�z�{a�  c3  �_݂�� *4  @� |  ɏ�����=��?��݆z���P  ) @@� h�݆z.�y��:���; ���� �z���`�z�' ꀁxzy�(2 	|�z��c6  b�  ��݂�_� :  ~0�| H�?� AՀ#K���9� ?}����������;��:��� c  ; ؐ��� by  :y �ȈB ����� 
  ~������z:�9�  ��  9�  ��0;  �>P�^���� ��A �� ��� �����: ߺ~��*�! ��� ���$�>;^&���cN  ; @@S9�{9 �:  �: :�� :U�Ҩ�bW  :�@@R��z� ��  �� :P9�� :/#��x����z' �@�x(9 	|�{Nsa�  b  �� :���:@ ?~I������� ";?��;W  ڸ�� c0  ;0 ـ��� cQ  ;Q ڈ�B ��b�  b�  c�  K��т^ʉ�Β^ϙ����z.���    ʡQ&��ݟ+Q��-� @�  :� �� ��� ��� ���ʚ��H  :@  �^ ��� �� ���ʚ�:?�`��<��>��  �� :q ӈ�bx  ;@@@SZ�{Z ;  ?)��S  �S 	�S 	B ���S �S :� ?~�����o����:_�`9���� bP  :P Ҁ��� a�  9� �p�B ����z8�;   �8  ;@  �^0:` �~P������� ��� ��� ��� �����:�ߺ}ߡ*� ��! ��>$�;>&���c8  ;@@@SZ�{Z �Y  �Y :� :��֘�b�  :�@@R��z� ��  �� 9�P:�� :4#�Ѡ�� �y�' �@�x(8 	|�{P�b  a�  � :��:� ?~������� ":���;S  ژ�� b�  :� �p�� cP  ;P ڀ�B ��8� bc  c�  K��т>ʊ�Β>Ϛ����z����    ��Q��`���m. @�  ;  �> �� ��{ ��ʚ~�H  :   �> ��� ��� ���ʚ��`   :�)`� �z�' ���x(. 	|�y��b  b�  ��:@ �^ ;@ �^+:� �:`@@Rs�zs �v  �v :   �>|:��:�:9���؈9�:����  ��  � �� � �� � �� �  �. "�  �/ "�+?) �A� ��[��[��^:�^>:`��~ �:������>�-� d@� p��0����*�*���v9�n~�q*: :; �9�:���;�����O  �X  �O �X �O �X �O �X �O  �o "�X  �x "��|��#H  @:   �>�:�  ��  :� ���:���b�  c�  H ������� ���. dA� \�>��> ��\ �9���;_� �~�� ����{Q' ���x(1 	|�z��b�  cU    �˓�ӫ.$�;,9�� "bd  a�  	�bB  N�!H  |��+C) �A� :  � H  d; Փ>:  �>  :� ���;_��cC  c�  H �)�)�z��:` �v  ��)����;  �  :@ �^�:��b  c�  H ��> )� �:  @� :   .1  A�	:�  �� �^ �) �:� A� :�  -�  A����z��:�  ��  9�  ��09� ��P���^��A �� �� ��! ��?��: ߺ~�*�� ��A ��^$��:�&���b�  :�@@Rրz� ��  �� :� 9��Ϙ�a�  :@@@RR�zR �O  �O ;P;?� :#��Ȉ� �{' ���x(: 	|�z�b4  c  �� :���:ݐ���zr' ���x(2 	|�y�sa�  by  � "b�  c�  H X��^ʊ�Γ^Ϛ����z5���  . @�  :@   ͇։�tm�cF�n�^ ��� ��{ ���ʚ~�H  9�  �� ��; �� ��>ʛ����z��:   �  :   �>0:�  ��P��^�A ��� ��� ��a Ȳ��9�ߺ}�q*�! �� ȳ$�>:�&���b�  : @@R�z �  � ;_� ::��Јb5  :@@@RR�zR �Q  �Q :�P:� 9�#�Ϙ����z�' � �x(8 	|�{.sa�  b�  �� :��b  c�  H Y`z  cU  ���^ʊ>Β^Ϛ>��^�zx��8  - @�  :� �� ��� ��� ���ʚ��H  :�  �� ��� �� ���ʚ��~�����_ݐH 0�> �)� �:@ A� :@  .2  A� :�`? M]c}%�  ;3 ٘�c4  9�@@Q΀y� :� ?~����  �� 	�� 	B ���� :� ?~�����o����:�`:����P   �s�9�_�J��b  : �Ј�U b�  :� Ո�B �����z��:�  ��  ;   �>09� ��P���>��! ��� ��A Тa ز��:@ߺ_�*�� Т� ز�$��:�&���b�  ; @@S9�{9 �4  �4 9�� :/��x�b.  :`@@Rs�zs �q  �q ;^P:_� :�#�א����{X' � �x(8 	|�{6�b�  cO  �� :���:` ?~i����� ":?��:T  Ҡ��� b:  :: �Ј�� bV  :V Ұ�B ��8� b�  c�  K��u��ʊ~Β�Ϛ~���{6��V  - @�  9� �� ��� ��� ���ʚ��H  :�  �� ��{ �� ��~ʛ�H �> �)� `:� A� :�  .6  A��;_�`>�M]b�}%��  : �Јb  : @@R1�z1 9� ?}���0  �0 	�0 	B ���0 9� ?  ϻ(��9^��}�����o����:��`:��� b�  :� Ԩ�� bz  :z �ЈB �����y��:   �2  :   �0:� ��P���^��A ��� �� �! �?��; ߺ~��*�� �� ��$��:>&���b2  : @@R�z �  � :�� ;W�ڸ�cV  ; @@S9�{9 �:  �: :�P;� 9�#�������z�' � �x(2 	|�zsa�  b�  � :���:� ?~������ ";_��:W  Ҹ�� cU  ;U ڨ�� bN  :N �p�B ��8� b�  c�  K��]��ʊ�Α�Ϛ����{.���  - @�  :  �> �� ��� ��ʚ��H  9�  �� ��� �� ���ʛ�;?�`=�M]a�}%��  :� �Ȉb�  :�@@R��z� :@ ?~I���  �� 	�� 	B ���� ;@ ?I���o  �i��� ]\������:��`9���� b�  :� װ�� a�  9� �p�B ���^�zt�:�  ��  ;@  �^0:  �>P������ �� ��� �! ��?��; ߺ~��*�A �a ��~$�^:�&���b�  ;@@@SZ�{Z �U  �U :?� 9��Έ�a�  ; @@S9�{9 �.  �. :�P;� :x#�����@�z�' �@�x(4 	|�{R�bT  b�  �� :?��:  ?~	����� "9���;Q  ڈ�� a�  9� ΰ��� cR  ;R ڐ�B ��8� b#  c�  K��e�~ʊΒ~Ϛ���{2���  -� @�  :� �� ��� ��; ���ʚ>�H  :`  �~ �� �� ��ʛ�;   �> :@  �^ AՀ#K��:�  �� ���y��;@  �W  :�  ��0:� ��P�>��~��a�! � �  �He�7 ������ճ��; ߺ~�*�A ����$�^9�&���a�  ;@@@SZ�{Z �N  �N :�� :��ո�b�  :`@@Rs�zs �u  �u :>P;� :#����� �z6' �@�x(6 	|�zY�c.  b/  �� ;_��:�ݐꀁz�' ꠁx(3 	|�z��b�  b�  � "cC  c�  H O��ʊ�ΓϚ����{2���  . @�  9� �� ��{ ��� ��~ʚ��H  :�  �� ��� ��; ���ʚ>�AՀ#K��X:   � `   ;^)`���{X' � �x(8 	|�{6�b�  cO  ���:@ �^+:~ �:�@@R��z� ��  �� :�  ��|:��: ::��؈;:����0  �8  �0 �8 �0 �8 �0 �8 �P  �� "�X  �� "9�  ���9� �� �\ �:���:~@�� �ꀁzq' � �x(1 	  ғ�$�`6]�T�Ğ|�{4�b�  bo  �� "8� �b�  ~��bB  N�!:��@�z' � �x(6 	|�{�cX  b  �)�� �z' ꀁx(3 	|�z��b.  b  ��)����� ����- dA� X�^��^ ��� �;_��;?� ���| �ꀁ{0' � �x(0 	|�z4�b�  c/  �� "c  cC  ~i�b�  N�!:�  �� H H:�� :W TҸ�bP  :   �2  �2 ;7 dٸ�c4  9�  ��  �� 9� yθ�a�  ;@  �N  :~@���zu' � �x(5 	|�z�b�  bq  ��B�[ ��(��ߖ9�ߎ~_y*;  
�?�p:�  ���0���8� �zz' ���x(: 	|�y��c  bu  ��ߢ:�ݠ: @@R1�z1 :  ~	��6  �6 	�6 	B ���6 :@  �_ݐ9�  ��ݔ;   �?ݖ:�  ��ݘ;_� 9�@@Q΀y�   ӈ���[l$�Ti�`:` ~i���  �� 	�� 	B ���� AՀ#K���AՀ#K���A݁�8!�� (|�����N� !        ����[�D��        �����������|�� (�!��`[  �A  < D� c�  ;�j�?� ��A݀�B (`|  �;  c>  �>�) A�  ;  �>�;=fp?9 c#  cb  H �H JH�>�)� A� H K@;  �>�;   �> �>(;  �|  �4���>(�(�  �>  .9�A� �  -8  A� ; ��>  �,
  ����  
  {  ��;��{  ��7�~��| H{d~�t��:��-�  z��~��@� ; ����7  ��;  6�|  �74Ȉ����  ��  .6�A� �>  -9  A� :����  �(4���>  
  {7  Ȉ  �� �H��RY��;��{  ��9�7�| Hz��tȈ;>%p-�  {7��@� :� ظ���  �>(c#  K��xw �b�  K��x� �� z���  ;=  :� �Ȉb�  �  �= �  �7 ?  =����z��� �z�' ꀁx{�(5 	|�z��b�  b�  �� �;   � 0�� 2. @� �>� ~��� �{4���  ) �@� h�� 2; ����� 0?  ~���� �z��:� ���� �z�����z�' ���xz��(8 	|�z��c6  b�  �� �AՀ#K��x� W6)� �@� h?  ~��� �z��z��;6��; ���ꀁ{5����{8' ꠁxzԣ(8 	|�z��b�  c3  �W �:� `��  � %c � %>� ~}��� ��� b:]  � f{5�~5��@� $z�' )4 	@�   �H[4Cὀ�g���zW' )� 	A� ��0Ր�~ҨP��0;  6�P|  �
  �= � �� @�� z�  ��:� @b�  b�  bE  K�3� 6�ٰ�� 2� | H�� @:�0�U  � �Y  � � @~��װ�� @2U | H�S @; ��8  �7  :�@ꠁz�' � �x(2 	|�{�b�  b�  � ��� @�� �] zU  ��b�  b�  b�  K�3�= �� �z��~X����bU  �� :� �6�| H{8  Ȉ:� @bC  b�  c  K�#:� ����z�' �@�x(9 	|�zV�b�  b�  � �:� ��� �] zV  ��b�  b�  b�  K�3�= �� �z��~�����b�  �� :� 6�| H{8  Ȉ:@ @b�  bD  c  K�#:� ?~��� ��r:� �֘�:�p՘�� b�  :� ֐�  �vT�#�*�J�� b�  :� ո�B �����z�' � �x(2 	|�{7�b�  b�  � �:@ ��] � *4  A� ��� ;  �| H>` ~]�� �z��~��װ�� �z��ꀁz�' � �xz��(5 	|�{�c4  b�  ����� )6  @� �>` ����z����  )� @@� p>� ~]����z��zx�;3��; ���ꠁ{4����{7' �`�xzի(7 	|�zu�b�  c7  ���� :� ~t�| H�} AՀ#K��p?  ~��:� ?~���U�U
r:�p֨�;
pب��V b�  :� ֠��X c  ; �ȈB ���� 
  ~�����^�zt�:�  ��  :@  �^0:` �~P������ x�� p�A p�a x�ub:�Z~U�*�� p�a x�~$��:^&���bT  :`@@Rs�zs   ���X���D�-��r  �r :�Pר�b�  :`@@Rs�zs �w  �w :^P:�fp>� ���`�zW' � �x(7 	|�z3�bp  bQ  � :�fp>� :@ ?~I��U
�W ":5
pѨ�:  и��Q b4  :4 Ѡ��P b  : Ш�B ��c$  b�  cb  K�w���ʊ�Β�Ϛ���^�zy���  . @�  :� �� ��� ��Z ���ʚ^�H  :`  �~ ��: ��� ��>ʚ��?  ~��: ��: ��� ��0  �� :� Ԁ�b�  :`@@Rs�zs ;  ?)��t  �t 	�t 	B ���t �t :� ?~��� ��r; �ذ�:�pհ��X c  ; �Ȉ�U b�  :� ՠ�B ����z7�:�  ��  ;   �>0:` �~P�^��� ��A ��! ��� ���b:�Z~6�*�! ��a ��~$�>:&  �%���oQUp���b  :�@@R��z� ��  �� :6PѰ�b7  :`@@Rs�zs �q  �q ;>P:]fp>R ��ꀁ{0' ���x(0 	|�z��b�  c1  � :}fp>s :� ?~���� ";6pٰ�:�  Ԙ��� c2  ;2 ِ��� b�  :� Ԉ�B ��8� bc  cb  K�u�ʊ>ΒϚ>����z���r  - @�  :  � ��: ��� ��>ʚ��H  :�  �� ��Z ��z ��^ʚ~�>� �:� ��:8�@� �4  :4 Ѡ�b6  :�@@R��z� :@ >~I���  �� 	�� 	B ���� �� :` ?~i�� ���r: ����;8p����� b  : А��� c1  ;1 و�B ���^�zu�:�  ��  :   �>0:� ��P���^��A ��� ��a ��� ���b:�Z~x�*  �ѓY9�߁T_ ؈�! ��� ���$�>:^&���bV  :�@@R��z� ��  �� :xP���bu  :�@@R��z� ��  �� :>P:�fp>� ��ꀁz2' ꠁx(2 	|�z��b�  b3  �V :�fp>� :� ?~���X�W ":8p���:�  Ը��Q b6  :6 Ѱ��T b�  :� Ԩ�B ��8� b�  cb  K�sՃʊ�ΓϚ���^�zv���  -� @�  ;  � ��� ��Z ���ʚ^�H  :`  �~ ��� ��� ���ʚ��?  ~�:� ��:H�P��T� �� �4  :T Ҡ�bS  :�@@Rրz� :� >~����  �� 	�� 	B ���� �� ;  ?)�� ���r; �؀�:0pр��X c  ; ظ��Q b6  :6 Ѱ�B ����z��:�  ��  :�  ��0:` �~P�^��  ڦ'QM���*wR�� ��A �� ��� ���b; Z~��*�� ��a ��~$��:�&���b�  :�@@Rրz� ��  �� :�PՀ�b�  :`@@Rs�zs �u  �u :�P:]fp>R �����z�' � �x(4 	|�{6��� :}fp>s :� ?~������ ":�pԀ�;3  ٘��� b�  :� Ԑ��� c5  ;5 ٨�B ��8� bc  cb  K�q��ʊ�ΒϚ�����z���r  . @�  :  � ��� ��� ���ʚ��H  :�  �� ��Z ��z ��^ʚ~�>  �;8 ��X�`��h�� ��  � :� �Ȉb�  :@@@RR�zR :` >~i��V  �V 	�V 	B ���V �V �V :  ?~)�� ���r: ����;8p����� b  : И��� c2  ;2 ِ�B ����z��:@  �Q    ��(���P���:`  �~0:� ��P������ ��� �� ��A ��Xb: Z~��*�a ��� ���$�~:�&���b�  :@@@RR�zR �T  �T :�P���b�  :�@@R��z� ��  �� :~P:�fp>� ���@�zt' � �x(4 	|�z2��V :�fp>� :� ?~���X�W ":�p���:7  Ѹ��T b�  :� ԰��Q b5  :5 Ѩ�B ��8� b�  cb  K�o��ʊ�ΓϚ���^�zv���  - @�  ;  � ��� ��Z ���ʚ^�H  :`  �~ ��� ��� ���ʚ�Ϋ>(:  ~9�|  �~44����(�(c  K��xu �b�  K��x� �] zS��}  :�  :� װ�b�  �=  �= �7  �7 >� �ꠁz��`�z' � �xzu�(6 	|�{5�b�  b    �2f.��)x�Hk�� �:   �= 0� 2-� @� �>@ ~}�� �{0���  * �@� h�� 2:� ~�����= 0>� ~]�� �{3�: И�ꠁz����z' ꀁxzի(1 	|�z��b�  b  � �AՀ#K��x�} Vw6) �@� h>� ~=�� �z��z�;��;9 �Ȉ�@�{����{' ꀁxz�(6 	|�z��bT  c  �� �:  `�  �= %c3 �} %>� ~ݺ� ��� �:]  � �z8�}���@� ${' *9 	@� zS' )3 	A� ��(ؐ�~��P��(:� ~��P|  �
  �� :  
� @::p;= @�q  �Q �Y �y  �� :� 
�Ȉ2� 
| H�� @z�  ��b�  c  b  K�3�6 @~Y��Ȉ�v @2� | H�� @:�\��  ��  � @~��Ȉ�6 @2q | H�v @  �b��K�zm��d~�:� ���  ��  :�@�@�z�' � �x(8 	|�z2�bP  b�  ���v @�} � z�  ��b�  c$  b�  K�3� ��z2�~r�Ӑ�bt  �= :� �~�| Hz  ��;  @bc  c  b%  K�#:V �ꀁzW' � �x(7 	|�{4�b�  bQ  ��:` ��} � {  ��bC  b�  b�  K�3�= ��z4�~t�Ӡ�bx  �] :� ~�| Hz  ��;  @bc  c$  b%  K�#:� ?~���V ��Vr; �ذ�:�pװ�� c  ; �Ȉ� b�  :� נ�B ���`�z�' ꀁx(2 	|�z��bp  b�  ��;  ��= �] )�  A� �� :� ~u�| H>  ~���{6�~V�Ұ����zT�ꠁzQ' � �xz��(1 	|�{�b�  bY  ��  ޖ:��c2�6w^�} *3  @� �>� ~����z5��U  ) @@� p>� =��Y�zx�{�:��:� а�ꀁz�ꠁz' �@�xz��(7 	|�zT�b�  b  �Y�� :� ~6�| H�= AՀ#K��p>� ~��:  ?~	��W�W"r:�pԸ�;7"pٸ�� b�  :� ���� c6  ;6 ٰ�B ��� 
  ~������z2�:�  ��  ;   �0:� ��P��>��! �� ��� ТA زWb; Z~��*� Т! ز>$��:&���b  :�@@Rրz� ��  �� ;Pظ�c  :�@@R��z� ��  �� :^P:�fp>� ��� �zQ' ꠁx(1 	|�z��b  bO  �� ;fp? :  ?~)���"�� ":�"pո�:X  ���� b�  :� հ�� bO  :O �x�  �z��sP�&LXB ��bd  c  cb  K�h���ʊ�Α�Ϛ�����y���6  -� @�  :  � ��z �� ��~ʛ�H  :�  �� ��� ��� ���ʙ��>� ~=�;1 ��� ԊZ ֲ�  �Y :� �Ȉb�  :`@@Rs�zs ;  ?	��u  �u 	�u 	B ���u �u :� ?~���� ���&r:� �ֈ�:�&pԈ�� b�  :� ֐�� b�  :� Ԁ�B ���^�zu�:�  ��  9�  ��09� ��P��>��! �� �� �A �Qb:`Z�*�� ࢡ 貾$��9�&���a�  ; @@S9�{9 �/  �/ :PЈ�b  ; @@S�{ �  � :~P:�fp>� �����zn' � �x(. 	|�{7�b�  bo  �� :]fp>R ;  ?	��&� ":&pЈ�:r  Ӑ��� b  :   ������-�#d�Cxи��� bu  :u Ө�B ��8� bC  cb  K�f��>ʋΓ>ϛ����y����  . @�  :� �� ��Z ��: ��^ʛ>�H  ;   � ��� ��� ���ʙ��>  ~��:� ���P�zT�V��  �t � :� נ�b�  ; @@S9�{9 ;  ?	��7  �7 	�7 	B ���7 9� ?}���� ���*r:5 �Ѩ�:�*p֨��Q b0  :0 р��V b�  :� ֠�B ����{7�9�  ��  9�  ��0:� ��P��~��a �� ��A � ��b; Z~U�*�� �� ���$��9�&���a�  :`@@Rs�zs �n  �n :PШ�b  :@@@RR�zR �P  �P ;>P:�fp>� �����{4' �`�x(4 	|�zo{a�  c3  �W 9�fp=� ;  ?	��*� ":*p  ��(EP����Ш�:�  �p��P b  : �x��T b�  :� Ը�B ��8� a�  cb  K�du�>ʋΓ>ϛ����y����  - @�  :` �~ ��Z ��: ��^ʛ>�H  ;   � ��� ��� ���ʙ�Ϊ�(��  ��  -��A� ��  .6  A� : ��>  ��,
  ~�����~  
  zr  ��;2��{8  Ȉ8��| Hy�d}�t��:��-/  z��~7z@� :� Ѱ��  ��(b�  K��xs �bc  K��x� �] zY��=  ;  :� ���b�  ��  �� ��  �� >� ~�� �y���`�y�' � �xzq�(2 	|�{1�b6  a�  ���;   � 0�� 2-� @� �>� ~���T�zy���  * �@� h�= 2:� ~������ 0>  ����y��:U   �#� ������Ҩ�ꀁzS�� �zQ' ���x{4�(1 	|�z��b�  bO  ���AՀ#K��x�� V�6) �@� h>� ~}���{1�z7�:Q��:� Ҹ�ꀁzO����zV' � �xyԣ(6 	|�z�b�  bY  ��:� `��  �= %b7 �� %=� }�z���:�  �Azp�}���@� $z' *4 	@� z�' )5 	A� �! а�~6�P�! :� }�P|  �
  �� �= �. @� {  ��:} @bc  b  bE  K�3� ~��՘��� 26 | H�. @:�0��  �7 ��  �5 � @~�И��N @2� | H�� @:� ��6  �0  :�@���z�' ꠁx(9 	|�z�{a�  b�  ��� @� �] zT  ��b�  bd  b�  K�3�� ��{5�}��Ϩ�a�  � :@ �~p�  �<1X�W���c^| Hzt  ��;  @a�  c  b�  K�#;. ����{5' � �x(5 	|�z6�b�  c3  �N�:  �� �� y�  x�c#  b�  c  K�3� ��z5�~բ֨�b�  �] 9� 2x| H{8  Ȉ:  @b�  b  c  K�#:  ?~)�� ���.r:n ��p�9�.p�p�� br  :r Ӑ�� a�  9� ϰ�B ��� �z�' ꠁx(1 	|�z��b  b�  ��:� ��� �� )�  A� ��] :  ~��| H>� ~���{.�~���p����z���`�z�' � �xzv�(2 	|�z6�b�  b�  ���� *7  @� �>� }ݪ�N�zo��/  ) @@� p>� ~ݢ��{0�z�:���:� ո��@�z���`�z�' � �xzr�(/ 	|�z2�bX  b�  ���   �-�Wz�D��Ҥ��:  ~�| H�� AՀ#K��p=� ~}r9� ?}���.�2r:�.p՘�:S2pҘ�� b�  :� հ�� bT  :T Ҡ�B ���� 
  ~������z/�:�  ��  :�  ��0;  �>P���������!�3b:�Z~�*������$��;>&���c7  ; @@S�{ �  � :3Pј�b0  :�@@R��z� ��  �� :�P9�fp=� �����z�' � �x(8 	|�{7�b�  b�  � :�fp>� ;  ?	��2� ":�2p֘�:�  נ�� b�  :� �x�� b�  :� �ȈB ��a�  b�  cb  K�]�ʊ~ΓϚ~���{/��/  -� @�  :  � ��� ��� ���ʚ��H  :`  �~ �� ��: ��ʛ>�=� ~=z:Q ��� �  �^�7�1p��c��@�� ���  �� :� ֐�b�  9�@@Q΀y� :� ?~����  �� 	�� 	B ���� �� :` ?~i�� ��6r9� �ψ�:�6pՈ��� a�  9� ϐ��� b�  :� Հ�B ���^�zt�9�  ��  ;   �>0;  �P������(� �� �A(�Qb:`Z~љ*�� ��(��$��;>&���c8  :�@@R��z� ��  �� :PЈ�b  :�@@Rրz� ��  �� :~P:�fp>� �����zx' ���x(8 	|�z�sa�  by  � :]fp>R :� ?~����6�� ":6pЈ�:r  Ӑ�� b  : �p�� bt  :t Ӡ�B ��8� bC  cb  K�[	��ʊ�Β�Ϛ����{1���  . @�  9� �� ��Z ��� ��^ʚ��H  :�  �� �� ��: ���  ��n)aaCGX�>Ϊ>(:� ~��|  �b�  K��`o  `�  a�  bd  K��`�  `�  `�  z  >� ~ݺ�� T�V \� P; p;8 ���c4  :6 P:� c#  b$  b�  K�3���z�����z�' �@�xz�{(. 	|�zO{a�  b�  ��:   � 0�= 2- @� �>� ~}����z���N  )� �@� h� 29� }��x��= 0?  ~���z��:� ֈ��`�z�����z�' ���xyӛ(2 	|�y�bx  b�  ��AՀ#K��x>� ~���5 cV76* �@� h=� ~]r���y��z��;6��:s ٘�� �{0�ꀁ{5' � �xz��(5 	|�z8�c  c7  ���9� `��  �� �a� �r �>  ~�����2:� p��6z��}8��@� ${' )� 	@� z�' *9 	A� ��ب�  �:G�壶
^����}��P��:` ~O�P|  �
  �] :  �4 @:�:� @��  ��  �� ;6 ٰ�2� | H�� @y�  p�c#  c  a�  K�3�t @~V�Ұ��4 @2 | H� @:�\��  ��  �� @6rٰ�� @1� | H�� @:z ��3  �9  :@���z' �@�x(5 	|�zW�b�  b  ���� @� �} zq  ��b  b�  b%  K�3�= ���z��~U�Ҩ�bO  �� ;  �~n�| Hzq  ��:� @bC  b�  b%  K�#:� �� �z�' ���x(5 	|�y��c2  b�  �T�;  �� �� y�  p�b�  b  b�  K�3�= ���y��5�٨�c3  �] ;  ~��| Hz�  ��9� @c#  a�  b�  K�#9� ?}���T ��T:r:4 �Ѡ�:�:pՠ��� b8  :8   �_��sg6ne�F3����� b�  :� �ȈB �����z' �`�x(/ 	|�znsa�  b  ��:@ ��] �� )7  A� ��� 9� ~o�| H>  }݂��{4�~T�Ҡ����zU�� �zV' ���xz7�(6 	|�y��b�  bY  ��� )�  @� �>` ~����z5���  * @@� p=� ~]z���z��{8�9���; ����`�y��ꀁy�' ꠁxz��(1 	|�z��bv  a�  ����� ;  x| H� AՀ#K��p>  ~��:  ?~)��T:�T>r:�:pՠ�9�>pΠ��� b�  :� �x��� a�  9� �ȈB ��� 
  ����^�zq�;   �1  9�  ��0:� ��P�����H��@�A@�aH�tb; Z~T�*�!@��H��$�>:�&���b�  :�@@Rր  ����}�z?���"z� ��  �� :tPӠ�br  ; @@S9�{9 �3  �3 9�P:=fp>1 ��� �y�' ���x(6 	|�z��c  a�  �Q ;=fp?9 :� ?~����>�� "9�>pϠ�;  �Ȉ�O a�  9� ψ��X c  ; ظ�B ��b  c#  cb  K�S���ʊ�Β�Ϛ�����z���q  - @�  :@ �^ �� ��: ��ʛ>�H  :�  �� ��� ��� ���ʚ��>  ~}�9� ��� ԋ ֲ�  � 9� �p�a�  : @@R�z ;  ?)��  � 	� 	B ��� � :� ?~���� ���Br:3 �ј�:�Bp՘�� b.  :. �p�� b�  :� Ր�B �����y��:�  ��  :�  ��0:� ��P�^�>��!X�AP�P��X��b9�Zy*�P�X�$��  ��R�"��tPt�g:�&���b�  ; @@S9�{9 �7  �7 :SPҘ�bN  ; @@S�{ �  � 9�P:fp> ��ꀁy�' � �x(6 	|�{4�b�  a�  �� 9�fp=� ;  ?	��B� ":SBpҘ�9�  �p��� bT  :T Ҡ��� a�  9� π�B ��8� a�  cb  K�Q�>ʋΓ>ϛ����z���  -� @�  :� �� ��� ��: ���ʛ>�H  ;   � ��� ��� ���ʚ��>` ~�:� ��:�����Z��5  �� �U :� Ԩ�b�  ; @@S9�{9 ;  ?	��4  �4 	�4 	B ���4 :� ?~���� ���Fr:p �Ӏ�:0Fpр��� br  :r Ӑ��� b5  :5 Ѩ�B ����{4�:�  ��  :�  ��0:� ��P�^�����h�A`��`�h�b  �o��T�6���; Z}��*��`��h��$��:�&���b�  9�@@Q�y� ��  �� :PPҀ�bX  9�@@Q΀y� ��  �� ;>P:�fp>� �����{5' ���x(5 	|�y��b�  c/  �� :�fp>� ;  ?	��F�� ":PFpҀ�;6  ٰ��� bW  :W Ҹ��� c8  ;8 ���B ��8� b�  cb  K�O͂�ʊ�Β�Ϛ�����z���  . @�  9� �� ��� ��� ���ʚ��H  :�  �� ��� ��� ���ʚ�΂,
  ~���>  ~}��0;3 ��Zl��n�Y  �� 9� �Ȉa�  :�@@R��z� :� ?~����  �� 	�� 	B ���� �� :� ?~��� ��Jr; �ؘ�:SJpҘ��� c  ; �Ȉ�� bU  :U Ҩ�B �����z��:   �4  :     � zbd�G�gq���0:� ��P�>�����x�!p��p��x��b:�Z}ӹ*�!p��x��$�>:&���b  9�@@Q�y� ��  �� ;3P٘�c6  9�@@Q΀y� ��  �� :�P:�fp>� ��� �z�' ���x(5 	|�y�b.  b�  �� :fp> :� ?~���J�� ";3Jp٘�:�  ׀��� c1  ;1 و��� b�  :� װ�B ��8� b  cb  K�M���ʊ�Β�Ϛ����z3���  - @�  9� �� ��� ��� ���ʚ��H  :�  �� �� ��: ��ʚ>Ϊ~bc  K��xv �b�  K��x� �] zX��  :�  ;7 ٸ�c/  ��  �� ��  �� >� ~�� �y�����y�' � �xzы(2 	|�{�b6  a�  ���9�  �� 0� 2-� @� �  �*�tD�_�F�ϲ#?  ~���T�zx���  * �@� h�= 2:� ~������ 0>  }݂��z��:Y �Ȉ�`�zX����zQ' ���xy�(1 	|�z�bt  bU  ���AՀ#K��x�� V�6) �@� h?  ����y��z7�:Q��:� Ҹ��`�zU�ꀁzV' � �xz��(6 	|�z�bn  bO  ���;  `�2  �= %b7 �� %>� ~���T��A�:�  ���y��}���@� $z' *8 	@� z�' )9 	A� �!а�~6�P�!:� ~��P|  �
  �� :` �t @:Z�9� @��  ��  � ;. �p�2� | H�� @{  ��c#  b  b%  K�3�� @~���p��t @2S | H�T @9����  � ��  � �4 @~��p��4 @2� | H�� @:z ��S  �P  9�@���y�'   �MO%?>�9;��ꠁx(8 	|�z��b�  a�  ���4 @�= �� z�  ��a�  a�  be  K�3�] ��{0�~��Հ�b�  �= :� �}Ѹ| Hy�  p�;  @b�  c  be  K�#;4 ��@�{0' ���x(0 	|�zғbV  c7  ���:  ��= �� y�  p�c#  a�  b�  K�3� �T�zp�~��׀�b�  �= 9� 1p| H{5  Ȉ:@ @b�  bD  b�  K�#:` ?~i�� ��Nr; �ؠ�:�Np֠��X c  ; �p��V b�  :� �ȈB �����y�' � �x(5 	|�z7�b�  a�  �T�:  �� �= )�  A� ��� :� ~5p| H=� ~�z�W�zt�~�Р�� �z�� �z' ꠁx{�(. 	|�z��c.  b  ����] *2  @� �>` ~=���  ��{�����@�Gz���  ) @@� p>  =����y��z��:w��:R Ӑ�ꀁzq�ꠁzv' � �xz��(6 	|�{�b�  bo  ���� :� ~W�| H�] AՀ#K��p>  ~��:� ?~���UN�URr;Npب�:�RpԨ��� c  ; �Ȉ�� b�  :� Ԁ�B ���� 
  ~�����^�zv�:   �  ;   �>09� ��P������������A��a��ub: Z~U�*����!��>$��9�&���a�  9�@@Q΀y� ��  �� :uPӨ�br  : @@R�z �  � ;>P:�fp>� �����{.' ���x(. 	|�y��b�  c3  �V :fp> 9� ?}����R�� ";5Rp٨�:�  ׀��Y c6  ;6 ٰ��W b�  :� �x�B ��b$  b  cb  K�F����  ��A�Q8��[q[��Α�Ϛ�����y���v  -� @�  :@ �^ ��: �� ��>ʚ�H  :�  �� ��� ��� ���ʙ�Ϊ� b�  K��xs �bc  K��x� �� z���  :�  ;7 ٸ�c2  �=  � �9  � >� }ݪ���zV��`�zT' � �xzo{(4 	|�{{a�  bW  ���:   �= 0� 2. @� �?  ~���U�zt��  ) �@� h�� 2:� ~������ 0=� ~=r��{0�:P Ҁ�ꠁzS�ꀁzO' ���xz��(/ 	|�z��b�  bY  ��AՀ#K��x�� V�6)� �@� h>  ~}����y��z��:T��:� Ҹ�ꠁzY�� �zQ' ���x{�(1 	|�zիb�  bO  ���:  `�  �� %b� �� %?  �����:�  ��z��~/��  �シDr2Ë��J@� $y�' ). 	@� z�' )� 	A� �Aϰ�~VxP�A:� 2�P|  �
  �= :  �8 @:�:� @�  ��  �� :t Ӡ�2� | H�� @y�  p�bc  a�  bE  K�3�� @4�٠��8 @2 | H� @:� ��  ��  ��$�~}�P|  �a�  K��`r  `�  bC  b�  K��`�  `�  `�  z�  �8 T� \�� P:� p:� ֨�b�  9� P:` b�  a�  be  K�3���{2����{1' � �xz�{(1 	|�z{a�  c5  ���:�  �� 0�� 2. @� �>` ~]����z���  ) �@� h�= 29� }��x��� 0>� ��X�zn�:� �p����z��� �z�' ���xz�(9 	|�y��b�  b�  ���AՀ#K��x>@ ~}��� cU�6)� �@� h>    �%��$��Wwh�=����y��z��:���:� ո�ꀁz���@�z�' � �xzT�(3 	|�z4�b�  b�  ���:  `�  �� �b� �� �?  ~]�����:r p���y��~4��@� $z�' )5 	@� zv' )� 	A� �� Ԙ�~�P�� ;  �P|  �
  � �= � @9� @}��p�� @~Ո| H�� @z3  ��a�  b�  be  K�3�� @.��p�� @2 | H� @:���  �5 ��  �9 �� @~�z�p��r @2� | H�� @; ��  �  :�@���z�' � �x(1 	|�{6�b�  b�  ��� @�� �} zw  ��b�  a�  b�  K�3� �z4�4�٠�c6  �� :` �}Ϙ| Hy�  p�:  @c#  b  b�  K�#:2 �� �z4' ���x(4 	|�z��  �;}Rs��C����c  b/  ��:` ��} �= {0  Ȉb#  b�  b  K�3�� ��y��~Ժ֠�b�  �} ;  ~3�| Hz0  ��9� @b�  a�  b  K�#9� ?}���� ���Vr:� �Ԑ�;Vpؐ�� b�  :� �Ȉ� c  ; ؘ�B �����z�' ���x(/ 	|�z�sa�  b�  �:� ��� �} *3  A� ��= 9� ~��| H>� }ݪ�z2�~Һ֐��`�z��ꀁz�' ���xz��(9 	|�y�bt  b�  ��� )0  @� �>  ~���{2���  )� @@� p>� ~}��z��y��:.��: р�� �z7�� �z2' ���x{8�(2 	|�y��c  b5  ���� 9� ~�| H� AՀ#K��p>� =�:@ ?~I���V��Zr:9Vp�Ȉ;Zp  �Ů��b���U����Ȉ� b3  :3 ј��� c  ; ذ�B ��� 
  ~������y��:�  ��  :`  �~0:� ��P�������������ȱ�b:�Z}ٱ*�A��aȲ~$�^:�&���b�  :�@@R��z� ��  �� 9�P�Ȉa�  :�@@Rրz� ��  �� :~P:]fp>R ��� �zt' ꠁx(4 	|�z��b  bo  �� :�fp>� :� ?~���Z�� ":yZp�Ȉ:  а��� br  :r Ӑ��� b  : Ш�B ��b�  b�  cb  K�=Y��ʋ>Β�ϛ>���z����  . @�  9� �� ��� ��� ���ʚ��H  ;   �> ��� ��� ���ʚ�Ϊ^&bC  K��xo �a�  K��x� � {��=  :  :p Ӏ�bn  ��  �� ��  ��   �޾\�K��c!0A�?  ~��ꠁy�����y�' � �xy��(8 	|�z5�b�  a�  ��:   � 0�} 2- @� �?  ~]���y���8  )� �@� h� 2:� ~������ 0>� ~��Pzy�9� �Ȉ���y��� �y�' ���xz/{(5 	|�z�{a�  a�  �PAՀ#K��x�� V�6* �@� h?  ��z5�z��9���:� θ����y���@�y�' ꀁxzO{(6 	|�z�{a�  a�  �;  `�.  �� %b� �� %>` ~]������:�  ��z4�}4��@� $z�' )� 	@� z�' *9 	A� ��԰�~��P���:� ~u�P|  �
  �} �� �� @�� y�  p�:= @b#  b�  b  K�3� 1�و��� 2� | H�� @:�L�w  �� �y  �� �� @~�r  ��L
9���\�Ԉ�� @3 | H� @:� ���  ��  :�@�`�z�' � �x(/ 	|�{3�bt  b�  ���� @�� � z  ��b�  b$  c  K�3�� ��y��~y��Ȉbu  � :  �~4�| Hz8  ��9� @bc  a�  c  K�#9� ����y�' ꠁx(9 	|�z��b�  a�  �:� ��� �} zn  ��a�  b�  a�  K�3� �z��~���Ȉb�  � :` }�| Hy�  x�:� @b�  b�  a�  K�#:� ?~��� ��^r:2 �ѐ�:r^pӐ��� b0  :0 р��� bv  :v Ӱ�B ��ꀁz�' � �x(5 	|�{4�b�  b�  ��;  �� �� )6  A� �� :� 5�| H>� ~����y���ؐ����{�� �{' ꠁxz6�(0 	  ��F�2�ҭx�
�6|�z��b�  c  ��"�� )�  @� �?  ~]��&z3���  * @@� p?  ~����&y��z��;4��:� ٸ�� �{2�� �{3' ꠁxz0�(3 	|�z��b  c/  ��"� :� ~��| H�� AՀ#K��p>@ ~=�:` ?~i��^��br;1^pو�:bpЈ��� c6  ;6 ٰ��� b  : ���B ���� 
  ~������z��;   �  :�  ��09� ��P������������ࢡ貱b; Z~��*�a����$�~9�&���a�  9�@@Q΀y� ��  �� :�PՈ�b�  ; @@S�{ �  � :�P:}fp>s �����z�' ���x(. 	|�y��b�  b�  �� ;fp? 9� ?}����b�� ":�bpֈ�:�  ���� b�  :�   ���YD$-+�7�֘��� b�  :� �x�B ��bD  c  cb  K�6���ʊ>Α�Ϛ>����y����  - @�  :� �� ��Z �� ��^ʛ�H  :   �> ��� ��� ���ʙ��>` ~���2~���c7  ���:� ��4H  :�  �� >@ ��84)� A� X�� �9�fp=� >` ~�;0��� �ꠁ{7' ꀁx(7 	|�z��b�  c1  � "8� �a�  ~��a�  N�!H >@ �:`  �x4:��:� TԸ�b�  :�  ��  �� :7 dѸ�b0  9�  ��  �� :� yָ�b�  :@  �V  :~@� �zu' ꀁx(5 	|�z��c.  bo  ������:��86:�.~�*:@ 
�X:�  ������ꠁzt' � �x(4 	|�{5�b�  bo  ��B:   �80:@:�@@R��z�   �Ì/�oD�<:��:@ ~I���  �� 	�� 	B ���� AՀ#K���AՀ#K������b�  A݁�8!�� (|�����N� !        ����[�D��                 �            �����������|�� (�!��`[  �A  < D� c�  ;�*@?� ��A݀�B (`|  �;  c>  �>�) A�  ;  �>�;=&?9 c#  cb  H ��H ܋>�)� A� H �;  �>�;   �> ?  =�; ���������  �� :� ���b�  ; @@S�{ :� ?~���  � 	� 	B ��� � :� ?~���� ���; ��Ȉ:��Ȉ� c  ; ذ��� b�  :� ט�B ���^�zv�:�  ��  :�  ��0:@ �^P�~���� h�a `�� `�� h��:@�~ّ*� `�a h�~$  �}{����z�����:�&���b�  :@@@RR�zR �T  �T :y��Ȉbu  :�@@Rրz� ��  �� :^P:�&>� ��ꠁzV' �`�x(6 	|�zu�b�  bQ  � :�&>� :` ?~i���� ":Y�Ȉ:6  Ѱ�� bP  :P Ҁ��� b3  :3 ј�B ��8� b�  cb  K�1�>ʊ~Γ>Ϛ~���z����  . @�  ;  �> ��z ��� ��~ʚ��H  :�  �� �� ��� ��ʚ�΂�,
  ~����>  ~]���;2 ��z������ �y  :� 
�Ȉb�  :�@@Rրz� :� >~����  �� 	�� 	B ���� �� �� :  ?~)�� ��
:� �Ԑ�:r
Ӑ��� b�  :� Ԁ��� bu  :u Ө�B ����z9�;   �  :�  ��0:� ��P���  �T��q|0��*��� x�� p�! p� x�; �~2�*� p�� x��$��:&���b  ; @@S�{ �  � :2�ѐ�b9  :�@@R��z� ��  �� :�P:�&>� ��� �z�' � �x(0 	|�{8�c  b�  � :�&>� ;  ?)��
� ":�
Ր�;  ظ�� b�  :� հ�� c  ; �ȈB ��8� 
b�  cb  K�/��^ʋ>Β^ϛ>���z6���  - @�  :@ �^ ��: �� ��>ʚ�H  :   �> ��� ��� ���ʚ��>` ~��; ���P�ZT�:V��  �X �8 : ���b  :�@@Rրz� :� ?~����  �� 	�� 	B ���� :` ?~i�� ��:� �ՠ�:TҠ�� b�  :� ո�� bV  :V Ұ�B ����{3�:�    �f��ξ�&�Ň���  :�  ��0:  �>P���� �� ��! ��� ���:`�4�*�� ��! ��>$��;&���c  :�@@Rրz� ��  �� ;4�٠�c3  : @@R1�z1 �9  �9 :�P:&> �����z�' �`�x(8 	|�zv��� :=&>1 ;  ?)����� ";ؠ�:q  ӈ��� c  ; ؀��� by  :y �ȈB ��8� b#  cb  K�-���ʋ>Β�ϛ>����z���0  -� @�  :� �� ��: ��� ��>ʚ��H  :�  �� �� ��: ��ʚ>Ϊ^(:� ~r�|  �~x4���(��(��  �>  .9�A� ��  -6  A� :����  �,
  ~����  
  z�  ��:r��zx  ��8��| Hz�d6t��:��-�  z��~��  �]�r�=�O%�R�@� : Հ��5  �^(bC  K��xs �bc  K��x� � {���  :�  ;4 ٠�c7  �  �= �  �9 >� ~]��`�z�����z�' � �xzӛ(4 	|�z�bp  b�  ��;   �= 0� 2. @� �?  ~���V�zt���  ) �@� h�= 2: ~����= 0>� ��X�zv�:� ԰����z��� �z�' ꠁxz�(9 	|�z��b�  b�  �X�AՀ#K��x�� V�6)� �@� h>  =���z��z��:W��:s Ҙ�� �zV�� �zP' ꀁxz8�(0 	|�z��c  bU  ���:� `��  �} %bv �� %>  ~����� �;  �� �z��~9��@� ${2' )2 	@� {' )� 	A� �! ����~8�P�! �:� ~��P|  �
  �� ��   �A�.B.��+�Q��� @�� z�  ��:} @bc  c$  bE  K�3� ~3�ј�� 2� | H�� @:�0��  �6 ��  �1 �P @�ؘ�� @2� | H�� @:� ���  ��  ;0�� �{2' ꠁx(2 	|�z��b6  c7  ���� @�� � {  ��c#  bd  bE  K�3� ���z��~��Ԉ�b�  �} :@ �~Ӑ| Hz�  ��:� @b�  b�  b�  K�#:0 �� �z2' �`�x(2 	|�zx�c  b5  ���:� ��� �� z�  ��b#  c$  bE  K�3�} ��z��~ؚ���b�  �= :@ ~��| Hz�  ��:` @b�  bd  b�  K�#;  ?	��� ���:P �Ҁ�:0р�� bS  :S Ҙ��� b8  :8 ���B �����{6' � �x(6 	|�{�b�  c5    �`ů��Т��ڃ����:` ��} �� *6  A� �� ;  ~��| H>� ~���T�zp�~кր�� �z��� �z�' �@�x{1�(5 	|�zQ�b2  b�  �T��� )7  @� �>  ���z����  )� @@� p>  ~}����z��zP�:���: Ԁ�� �z��� �z�' ���x{8�(1 	|�z��c  b�  ����] :  ~��| H�� AՀ#K��p?  ~=�:� ?~������;؈�:qӈ�� c  ; ؐ��� bp  :p Ӏ�B ���= 
  7�Ȉ��z��:   �  :@  �^0;  �>P����� ��� �� ��� ���:@�~�*�! ��� ���$�>:�&���b�  : @@R�z �  � :Q�҈�bU  ; @@S9�{9 �2  �2 :�P:&>    �Y�l��w���ꀁz�' � �x(5 	|�{4�b�  b�  �� :]&>R :� ?~������ ";1و�:�  ֐�� c0  ;0 ـ��� b�  :� �x�B ��b�  bC  cb  K�&1��ʊ>Α�Ϛ>����y����  . @�  :� �� ��� ��Z ���ʚ^�H  :   �> ��� ��� ���ʙ��� &z���p ?  ~���6�~��P|  �b�  K��`r  `�  bC  b$  K��`�  `�  `�  y�  �� T�� \�� P:� p: Ш�b  :v P;  b  bd  c%  K�3���{�� �{' ꀁxz7�(/ 	|�z��b�  c  ���9�  �� 0� 2- @� �>` =���z2���  )� �@� h� 2:� ~������ 0>� ~ݢ�V�zn�: �p�� �z����z' ���xy��  t "JI�jR#�J(8 	|�z��c4  b  ���AՀ#K��x>@ ~}��� cU�6* �@� h=� z���z��z�:���;9 �Ȉꀁz���`�z�' � �xzt�(. 	|�z4�b�  b�  ���:� `��  �� �b� � �?  ~]���� �:r p�� �y��}4��@� $z�' )� 	@� zu' *5 	A� �� �Ԙ�~�P�� �;  7�P|  �
  �= �= �2 @� z  ��9� @a�  b�  a�  K�3�� ~���x��} 2� | H�� @; ��8  �5  :2�� �z4' ���x(4 	|�yЃb  b7  ����r @�} � {  ��b#  a�  c%  K�3� ���z��}ԪΠ�a�  �} ;  �}��| Hy�  x�:� @a�  b�  c%  K�#:� �ꠁz�' � �x(4 	|�z�b�  b�    �!_�G/�5�2���;  �� �} zv  ��b�  b$  b�  K�3�= ��z��}��π�a�  � :` ~��| Hz�  ��:� @a�  b�  b�  K�#:� ?~��� ��: �А�9�ΐ��� b  : И��� a�  9� �x�B ��ꀁz5' � �x(5 	|�{4�b�  b7  ���;  �� �� )/  A� ��} :� 5�| H>  ~�����z���ؐ����{�� �{' ꠁxz{(3 	|�z�{a�  c  ���� )�  @� �>� =��Y�zn���  * @@� p?  }����z4�z��:���:� װ��@�z���`�z�' ꠁxzr�(. 	|�z��bP  b�  ��� :� ~��| H�� AՀ#K��p?  ~}�9� ?}�����:�ט�:SҘ��   �*ƍ�)'rQȂb�  :� �x�� bX  :X ���B ���� 
  ~������z��;   �  9�  ��0:  �>P������ �� �� ��� Ȳ�; �~��*�� ��� ȱ�$��:>&���b6  : @@R�z �  � :��՘�b�  ; @@S�{ �  � 9�P9�&=� �����y�' � �x(0 	|�z6�b�  a�  �� ;&? :  ?~	��� "9�Ϙ�:�  ���� a�  9� �p��� b�  :� ֈ�B ��c$  c  cb  K�a�ʊ~ΒϚ~���z.���  - @�  :� �� ��: �� ��>ʛ�H  :`  �~ �� ��: ��ʚ>�=� ~�r:U ���P��T��V��  �� �� :� Ԑ�b�  ; @@S�{ :` ?~i��  � 	� 	B ��  ��I*������ :  ?~	�� ��"9� �Ψ�:�"ר�� a�  9� ΰ�� b�  :� �x�B ���^�zt�:   �4  :   �09� ��P���>��! ��� �� ТA زU:`��*�! Т� ز�$�>:&���b  ; @@S9�{9 �0  �0 :��֨�b�  ; @@S�{ �  � :~P:�&>� ��� �zo' � �x(/ 	|�{1�b8  by  � :&> :@ ?~I��U"�P ":�"֨�9�  π�� b�  :� ֈ�� a�  9� Ϡ�B ��8� b  cb  K�I�~ʊ^Β~Ϛ^���z���1  -� @�  ;  � �� ��z ��ʚ~�H  :@  �^ ��� ��� ���ʚ��:   �> H ?  ~��9�`9� T�p�a�  ;   �  � : d�p�b    <^uK�.�H�0\�:@  �P  �P :� y�p�b�  :   �4  ;>@���{8' ���x(8 	|�y��b�  c3  �W���������:��~�*:  
�7�:�  ��p��x� �{/' ���x(/ 	|�z����:w�:@@@RR�zR 9� }���S  �S 	�S 	B ���S :   ��AՀ#K��4AՀ#K��<A݁�8!@� (|�����N� !    ����[�D�        �����������|�� (�!�A`[  �A  < D� c�  ;�B@?� ��A݀�B (`|  �;  c>  �>�) A�  ;  �>�;=>?9 c#  cb  H �H )ċ>�)� A� H *�;  �>�;   �> �>,
  8�Ȉ;>�:� �Ȉ�  ?  �:� P? �@c9�@{9�g9��c9�%�7  ;7 ٸ�c7  :�@@R��z� :� ?~����    ��T�.�Y�,�%�� 	�� 	B ��:� ?~���� _��;8 P���:����� c6  ;6 ٰ��� b�  :� ט�B ���^�zv�:�  ��  :�  ��0:@ �^P�~���� h�a `�� `�� h��:@�~ؑ*� `�a h�~$��:�&���b�  :@@@RR�zR �T  �T :x����bu  :�@@Rրz� ��  �� :^P:�>>� ��ꠁzV' �`�x(6 	|�zu�b�  bQ  � :�>>� :` ?~i���� ":X���:6  Ѱ�� bP  :P Ҁ��� b3  :3 ј�B ��8� b�  cb  K�A�ʊ~ΓϚ~���z����  . @�  ;  � ��z ��� ��~ʚ��H  :�  �� �� ��� ��ʚ��>� =�:9 P�Z �� ��Q  � :q ӈ�bt  :�@@R��z�   ��g޶��ͼ��:  ?~	���  �� 	�� 	B ���� �� :� ?~���� _��
:Y P�Ȉ;
�Ȉ� bT  :T Ҡ�� c  ; ب�B �����z��:�  ��  :�  ��0:  �>P������ x� p�� p�� x��:`�~��*� p�! x�>$��:�&���b�  :�@@R��z� ��  �� :���Ȉb�  : @@R1�z1 �7  �7 :�P:>> ��ꠁz�' �`�x(6 	|�zu�b�  b�  �� :=>>1 :` ?~i��
�� ":�
�Ȉ:�  ֈ�� b�  :� ׀��� b�  :� ֘�B ��8� b#  cb  K�-�>ʊ~Γ>Ϛ~���z���0  - @�  ;  �> ��z ��� ��~ʚ��H  :�  �� �� ��: ��ʚ>�?  ~]�:� P��ȃ:Њzԓ6 �v   �J{�		���al��  :� ԰�b�  : @@R�z :  >~)��  � 	� 	B ��� � � ;  ?	�� _�:r PӐ�:�א�� bv  :v Ӱ��� b�  :� ׈�B ����{0�:   �0  :�  ��0:� ��P���� ��� ��! ��! ��2: �2�*�� ��� ���$��;&���c  : @@R1�z1 �8  �8 ;2�ِ�c0  :�@@R��z� ��  �� :�P:�>>� ��� �z�' � �x(8 	|�z�b8  b�  � :�>>� :  ?~	��� ":�֐�;5  ٨�� b�  :� ���� c4  ;4 ٠�B ��8� b�  cb  K��^ʊ�Β^Ϛ����z8���  -� @�  :@ �^ ��� �� ���ʚ�H  :   �> �� ��� ��ʚ��  	�'�\�42�|p��b�  K��xs �bc  K��x� �= {6���  :]  :� Ԑ�b�  �=  � �4  � >� ~���`�z����z' � �xzӛ(2 	|�z3�bt  b  ��R;   � 0�= 2. @� �>� ~]��Vz3���  ) �@� h� 2:� ~����� 0?  ~���Vz2�:r Ӑ�ꠁzt����zx' � �xz��(8 	|�{5�b�  bq  �RAՀ#K��x�] VT6)� �@� h>� ��XVzy�{5�:9��:� Ѩ�� �z6�ꀁz7' �@�xz��(7 	|�zP�b  b3  �XR;  `�1  �� %b� �� %>� ~���W_�A �:  � �{1�~1��@� $z5' )5 	@� z' )� 	A� �xр�~��P��x:` ~T�P|  �
  �] ;  � @;:�:� @��    
4�G�T���q�O� �� ��  � �� �} :U Ҩ�3 | H� @zy  ��bC  b$  c%  K�3�� @~�Ш�� @3 | H� @:z ��S  �P  :7�� �z6' ꀁx(6 	|�z��c2  b3  �Wb� @� � z  ��b#  b�  b�  K�3� �f{3�~S�Ҙ�bP  � :� ��| H{  ��:� @bC  b�  c%  K�#:w P� �zv' ꠁx(6 	|�z��b  by  �b:@ ��] � z�  ��bc  b$  b�  K�3� �f{0�~P�Ҁ�bT  �} :� �| H{  ��:� @bC  b�  c%  K�#:  ?~	��W _�W:� PԸ�:�ָ�� b�  :� Ԩ�� b�  :� ր�B ���`�z2' � �x(2 	|�z�bx  b9  �b:� ��� �]   ��}��a����:*2  A� �� :  ~q�| H?  ���fz��~U�Ҩ�ꀁzP�� �zY' ���xz4�(9 	|�zԣb�  bW  ��r�} )3  @� �>� ~��v{1��Q  )� @@� p>� ~���Wvzv�z��;��:� ب�� �{�� �{' �@�xz0�(4 	|�zP�b  c  �Wr�� :� 5�| H�= AՀ#K��p>  ~��;  ?	��T�T:Р�:�נ�� b  : а�� b�  :� ר�B ���= 
  ~3�����{2�:�  ��  :�  ��0:  �>P��>��! �� �� ��A ��T:��~��*�! ��! ��>$�>;&���c  :�@@R��z� ��  �� :��֠�b�  : @@R1�z1 �6  �6 :^P:�>>� ��� �zY' � �x  긤���F�'�(9 	|�z8�c  bO  �� :�>>� ;  ?)����� ":4Ѡ�:V  Ұ�� b8  :8 ����� bY  :Y �ȈB ��bd  b�  cb  K�A��ʉ�Α�ϙ����{5���  . @�  :` �~ ��� ��� ���ʙ��H  9�  �� �� ��: ��ʛ>Ϊ�b�  K��xt �b�  K��x� �� z���  :]  :2 ѐ�b3  ��  �� ��  �� =� r� �zu�ꀁzw' � �xz��(7 	|�z�c.  bo  ��b:@  �] 0�� 2- @� �>  ~����fz���  )� �@� h�} 2;3 /�Ȉ�� 0=� r�fz2�:� ֐�ꠁz��ꀁz�' � �xz��(3 	|�{5�b�  b�  ��bAՀ#K��x� V6* �@� h>@ ~���Wf  <p���k.�8�zt�z��:���;9 �Ȉꠁz�����z�' � �xyի(8 	|�z�b�  b�  �b:@ `�V  �} %bt � %?  }���o�� �9�  � �z8�}8p�@� ${' )� 	@� y�' *2 	A� ��p�p�~��P��p:` 6�P|  �
  �= :� �� @:��: @~�xr7 A� �T  �� �P  �� H  �T �P �= :� Հ�29 | H�/ @{7  Ȉb�  c  b�  K�3�� @~��Ԁ��o @2S | H�O @:: �1  �4  ��b�  K��xx �c  K��x� �� z����  : �p�b  �]  �= �P  �0 � �zt�ꠁzx' ���xz��(8 	|�z��c0  bq  �r:�  �� 0�� 2- @� �>@ ~����vz���  )� �@� h�} 2;3 1�Ȉ  2PB^�2��Z�= 0>  }����vz��:N �p�ꀁzU�� �zS' � �x{�(3 	|�{4�b�  bQ  �rAՀ#K��x�� V�6* �@� h=� ~�r�Uvzx�{�:���;9 �Ȉ� �z�����z�' ���xy�(6 	|�z�b2  b�  �Ur9� `��  � %c �= %>  }������ �:=  �A �zu�}5��@� $z�' )� 	@� z4' *4 	A� �hՈ��P�h;  ~�P|  �
  � �� �� @:] @~r�Ӑ��� @~��| H�� @z�  ��bc  b�  b%  K�3� @2�ِ�� @2� | H�� @9� ���  ��  �� @~r�Ӑ�� @25 | H�/ @; ��  �  :�����z�' � �x(4 	|�{.sa�  b�  ����� @�� �= z8  ��b�  bD  c  K�3  (���X{c�� �O�zy�}ق�Ȉa�  � :� �~4�| Hz8  ��:@ @a�  bD  c  K�#:o P� �zy' ꠁx(9 	|�z��b  by  ��:� ��� � z�  ��bc  b�  b%  K�3�� ��z��~rА�b  � :� ~x�| Hzq  ��:� @b  b�  b%  K�#:� ?~��� _�9� P�x�:O�x�� a�  9� θ�� bS  :S Ҙ�B ��ꀁz�' � �x(5 	|�{4�b�  b�  ��;  �� �} )3  A� ��� :� 5�| H>� ~����z/���x��`�{����{' ꠁxyӛ(7 	|�z��bp  c  ���� )�  @� �?  }�����z����  * @@� p>� ��X�zq�z0�:���: Ԁ�� �z�����z�'   �6	,�7���,s���xy��(7 	|�y��c2  b�  �X�� :  ~�| H� AՀ#K��p>� }��:� ?~����9��x�:��x��N a�  9� Ψ��T b�  :� Ԉ�B ��� 
  ~�����{7�:   �7  :�  ��0:` �~P�^��� ��A �� У! س/: ��*�� Т� ز�$��:~&���bp  :@@@RR�zR �S  �S ;/��x�c8  : @@R1�z1 �9  �9 :�P:�>>� ��� �z�' �`�x(2 	|�zp�b  b�  � :=>>1 :@ ?~I��O�Q ":��x�:  Ј�� b�  :� ո�� b  : И�B ��b�  b#  cb  K���^ʉ�Β^ϙ���^�zw��7  - @�  ;  � ��� ��: ���ʚ>�H  9�    ,���~P��'A�� ��Z ��z ��^ʚ~�>� =�:� P�������  � �� ; ؠ�c  : @@R1�z1 9� ?}���8  �8 	�8 	B ���8 :@ ?~I��Y _�Y":� P�Ȉ9�"�Ȉ� b�  :� ׀��� a�  9� ΰ�B ����z/�;   �  :`  �~0:@ �^P������ ��� �� � �: �~��*� �� ��$�:~&���br  :�@@R��z� ��  �� :���Ȉb�  :�@@R��z� ��  �� :>P9�>=� ��� �z2' ꠁx(2 	|�z��c  b3  �O :>> :� ?~���"�� ":�"�Ȉ:0  р��V b�  :� ����Q b/  :/ �x�B ��8� b  cb  K�Ⴞʊ�Β�Ϛ����{/��o  -� @�  :@ �^ �  ߩ3E�8��� ��� ��ʚ��H  :�  �� �� ��: ��ʛ>�=� ~}z9�����(|�b�  a�  ��>� ~]�:��ꀁz�' � �x(8 	|�{4����AՀ#���| Ha�  �:� �w  ��~i�N� >� ���z��9� ��  ��>@ ~����z3���  ~6p A�
H  lH  h>� �:����(|�a�  b�  ���AՀ#K��L?  ~]���� ��A �zn���  :� }��|  �}�4x���  AՀ#K��x>� ��8�> ffb1fg> ffbffz ~QȒ~Rt{1�~R�R 
~R�P-2  :` A� :`  -�  A�>� ~��9� P:� %��  9� �x�a�  ; @@S�{ :  ?~	��  � 	� 	B ��� � � :  ?~)�� _�&:T PҠ�:t&Ӡ�  &1/����D��� bU  :U Ҩ��� bo  :o �x�B ����z.�;   �.  ;   �09� ��P�������� �� ��: �~ԉ*�! ����$�>;&���c  :�@@R��z� ��  �� :��ՠ�b�  :�@@Rրz� ��  �� :>P9�>=� ��� �z/' ���x(/ 	|�z��c6  b7  �� ;>? :  ?~	���&�� ":�&ՠ�:8  ����� b�  :� �Ȉ�� b0  :0 р�B ��8� c  cb  K��m��ʉ�Α�ϙ����{4��  . @�  :� �� ��� ��� ���ʙ��H  9�  �� �� ��: ��ʛ>�:�  �� >  ~}��S��^  �>  -1�A� �  -�  A� :����  ��  
  z�  ��9���y�  p�8��| H  �b�%���!5n��{4�~�t��:~%p.4  zr�~3�@� :R ѐ���  b�  K��xw �b�  K��x� �� z����  9�  ; �p�c  �=  �� �8  �� >` ~]�� �z����z' ���xz�(6 	|�y�b8  b  ��9�  �� 0� 2- @� �>` ~�����z���  )� �@� h�= 2;1 8�Ȉ� 0>@ }ݒ�N�zt�:� ֠�ꠁz�����z�' � �xy��(0 	|�z5�b�  b�  ��AՀ#K��x�] VS6* �@� h>� ~�����y��z�:���:1 ֈ�ꠁz��� �z�' �`�x{�(2 	|�zu�b�  b�  ���:� `��  � %b �= %?  ��X��A:�  ��y��}7��@� $z�' )� 	@� z�' *6 	A� �`ר�~�P�`  �)� ��Gˈ�F�:  0�P|  �
  �= :` �x @:Z 9� @��  ��  � :� �p�2� | H�� @z�  ��b�  b�  b  K�3�8 @.��p��x @2S | H�X @9�\��  ��  :�����z�' � �x(7 	|�z�b�  b�  ���x @�} �] zO  ��b�  a�  a�  K�3� ���z��~9��Ȉb0  �} :@ �}Ӑ| Hy�  p�:� @b#  b�  a�  K�#:� Pꠁz�' � �x(9 	|�z�b�  b�  �X�9� ��� �= z6  ��b�  b�  b�  K�3�� �X�zy�~z�Ȉb  �� :  ~�| Hz�  ��:@ @b  bD  b�  K�#:` ?~i��� _��*;8 P���:�*���� c7  ;7 ٸ�� b�  :� Ր�B �����z�' ���x(3 	|�y��  [+�ΗO���{bb�  b�  ��9� ��� �] )2  A� ��� :` }�| H>� ~ݢ��z8�}�z����@�y��� �y�' �`�x{2�(7 	|�zr�bP  a�  ��� )�  @� �=� z��z����  * @@� p>` }ݚ��z2�zV�9���:� ϰ�ꀁy��ꠁy�' ���xz��(9 	|�z��b�  a�  �N�� :  ~р| H�� AՀ#K��p?  ~��;  ?)���*��.9�*Ϩ�:�.Ԩ��O a�  9� �p��T b�  :� Ԁ�B ���= 
  ~8������z��:   �  9�  ��0:` �~P�^�>��!(�A �� ��(��: �~Ձ*�! ��(��$�>:~&���bq  :@@@RR�zR �S  �S :��ר�b�  : @@R�z �  � 9�P  ������2O(;=>?9 ��� �y�' �`�x(2 	|�zq�b6  a�  �� :>> :@ ?~I��U.�P "9�.Ψ�:0  р��� a�  9� �Ȉ�� b3  :3 ј�B ��c  b  cb  K��)�^ʊ�Β^Ϛ���^�zy���  - @�  :� �� �� �� ��ʚ�H  :�  �� ��Z ��z ��^ʚ~�AՀ#K���?  ~��:� P����:���  �4 9� Π�a�  ; @@S�{ :  ?~	��  � 	� 	B ��� � :� ?~���W _�W2;7 Pٸ�9�2ϸ�� c4  ;4 ٠�� a�  9� ϰ�B ����z��9�  ��  :`  �~0:@ �^P���>��!8��0�0��8��:��~�*��0�8�$��:~&���br  : @@R1�z1 �3  �3 :��ָ�  <"��a�_�g%U�b�  : @@R�z �  � :�P;>? �����z�' � �x(2 	|�z.sa�  b�  �X :�>>� :  ?~	��2� ":�2ָ�:�  ՠ��V b�  :� �p��U b�  :� ���B ��8� b�  cb  K���>ʊΒ>Ϛ��^�zw��  -� @�  9� �� ��� ��: ���ʚ>�H  :   � ��Z ��z ��^ʚ~�>� �9� P�: Ԋ� ֳ/  �� :� �x�b�  :�@@R��z� :  ?~)���  �� 	�� 	B ���� �� :  ?~	��X _�X6:� P���;86���� b�  :� �x��� c.  ;. �p�B ����z6�:`  �v  :@  �^09� ��P������H��@�@�H�: �~��*�a@��H��$�~:^&���bN  :�@@R��  �h���^��kz� ��  �� 9�����a�  :�@@R��z� ��  �� :>P:�>>� ���`�z.' ꠁx(. 	|�z��bn  b/  �� :]>>R :  ?~	��6�� ":86���:r  Ӑ��� b6  :6 Ѱ��� bp  :p Ӏ�B ��8� bC  cb  K�����ʊ�Β�Ϛ�����y���  . @�  :� �� ��Z ��� ��^ʚ��H  :�  �� ��� ��� ���ʙ��?  ~�;0 P��P�zT�:V��  �y �9 :� �Ȉb�  :�@@R��z� :� ?~����  �� 	�� 	B ���� 9� ?}���� _��:; P؀�:�:׀��X c  ; ؈��W b�  :� �ȈB ����z��9�  ��  9�  ��0;  �>P�>�~��aX�!P�AP��X��:��~P�*��P��X��$  jXnb�Җ��|t��9�&���a�  :`@@Rs�zs �n  �n :0�р�b4  :@@@RR�zR �Q  �Q :�P:�>>� �����z�' �`�x(9 	|�zo{a�  b�  �V 9�>=� :� ?~���:�� ":0:р�;.  �p��Q b/  :/ �x��Y c6  ;6 ٰ�B ��8� a�  cb  K��Ⴞʊ�Β�Ϛ�����y����  - @�  :` �~ ��Z ��� ��^ʚ��H  :�  �� ��� ��� ���ʙ��:   � H L>� ~��;`;8 T���c1  :`  �y  �y :X d���bU  :�  ��  �� 9� y���a�  :   �  :�@� �z�' � �x(3 	|�{1�b4  b�  ����Z �(��9��~Wy*�0��8�z<��زw���;7�� �{5' ꀁx(5 	|�z��b.  c/    �ˢ���o������b;  ��:@  �Wp�Wx�`�z�' ꠁx(0 	|�z��bx  b�  ��:�  ���:7�9�@@Q�y� 9� }����  �� 	�� 	B ���� AՀ#K��AՀ#K��A݁�8!�� (|�����N� !    ����[�D�        �����������|�� (�!��`[  �A  < D� c�  ;�&@?� ��A݀�B (`|  �;  c>  �>�) A�  ;  �>�;=" ?9 c#  cb  H _aH <�>�)� A� H $;  �>�;   �> �>,
  8�Ȉ�0?  �;8 ���@��D��  �� :� �Ȉb�  ; @@S9�{9 :� ?~���7  �7 	�7 	B ���7 �7 
:� ?~���� ���;8 ����:� ���� c6  ;6 ٰ��� b�  :� ט�B ���^�zv�:�    DlQ��P@�;�B��  :�  ��0:@ �^P�~���� h�a `�� `�� h���:@�~ؑ*� `�a h�~$��:�&���b�  :@@@RR�zR �T  �T :x����bu  :�@@Rրz� ��  �� :^P:�" >� ��ꠁzV' �`�x(6 	|�zu�b�  bQ  � :�" >� :` ?~i���� ":X ���:6  Ѱ�� bP  :P Ҁ��� b3  :3 ј�B ��8� b�  cb  K�흃ʊ~ΓϚ~���z����  . @�  ;  � ��z ��� ��~ʚ��H  :�  �� �� ��� ��ʚ�Ϊ�(;  ~7�|  �b#  K��`r  `�  bC  c  K��`�  `�  `�  zs  �� �� �}  : 0:� ր�b�  :� b�  c�  b�  K�3>  ~]�� �{4�ꠁ{3' � �xz��(3 	  x?��Re5�p�|�z���:�  �� P�� R- @� �>  ~���T�zu��  )� �@� h�= R; ����� P>� ~=��Q�zt�:� ՠ�� �z��� �z�' ���x{�(6 	|�z��b  b�  �Q�AՀ#K��x�� V�6* �@� h?  ~����z��z��:w��: Ӏ��@�zq�� �zx' ꀁx{2�(8 	|�z��bT  bu  ���:� `��  � Db �= D?  ����� r:] 0�� vz��}3��@� $zp' )� 	@� zQ' *1 	A� �! �Ӑ�2�P�! �:� ~��P|  �
  ��  :� �� `:� �: `�7  �0  �]  ;0 ـ�2� | H�� `zT  ��c#  bd  b�  K�3�� `~�׀��8 `2� | H�� `:Z ��2  �7  :x�ꀁzv' � �x(6 	|�z4�  -�욫_n[3�b�  bw  ���� `��  �]  zY  ��bc  b  c%  K�3�=  ���z��~��ՠ�b�  �  ;  �~��| Hz�  ��:  @b�  b$  b�  K�#:� ��@�z�' � �x(9 	|�z�bP  b�  ��:� ���  �  z�  ��b�  bd  b�  K�3�=  ��z2�~��֐�b�  �  :� ~�| Hz  ��;  @b�  c$  b%  K�#:@ ?~I�� ���
:� ����:
 ���� b�  :� װ��� b  : �ȈB ��� �zr' � �x(2 	|�{1�b4  bu  ���:� ���  �]  )2  A� ��=  :` ~3�| H>� ~�����z��~X����� �zY��`�zU' ���xzp�(5 	|�zЃb  bW  ����=  )�  @� �?  =��Y�zu��  * @@� p  c�W��5�d��k>� ~ݺ��z4�z��:T��; ���� �zS�ꠁzW' � �xz��(7 	|�z�c0  bQ  ���  ;  ~x�| H�}  AՀ#K��p>� ~��:@ ?~I��
�:7
 Ѹ�: и��Q b6  :6 Ѱ��P b  : Р�B ���  
  ~�����^�zx�:�  ��  :�  ��0:� ��P�^�~��a ��A �� �� ���:��~��*� ��a ��~$��:^&���bX  :�@@R��z� ��  �� :��ָ�b�  :�@@R��z� ��  �� ;P:�" >� ���@�{' ꠁx(3 	|�z��bN  c  �� :�" >� :` ?~i���� "; ظ�:V  Ұ��� c  ; ؘ��� bU  :U Ҩ�B ��c$  b�  cb  K��ɂ�ʊ�Β�Ϛ����   6��c9Xv�Ѓz����  - @�  9� �� ��: ��� ��>ʚ��H  :�  �� ��� ��� ���ʚ��>` }��:��:H�ZP�X� �0  �P 9� ΀�a�  :�@@Rրz� :� ~����  �� 	�� 	B ���� :� �ꠁz�' � �x(3 	|�{�b�  b�  ��:  ��=  �]  zW  ��b�  b  b�  K�3��  �O�zn�~���p�b�  �  :  ~��| Hz�  ��:@ @b�  bD  b�  K�#:` ?~i�� ��:� ��x�9� �x�� b�  :� ֈ��� a�  9� ΐ�B �����z' � �x(3 	|�{7�b�  b  ���;  ��  �]  )�  A� ��=  :` 3�| H>  ~����z����x��@�{����{' �`�xzғ(1 	|�zr�bT  c  ���  ! �i��.*ӡp��  *0  @� �?  }����z.���  ) @@� p>` ���z��zW�;2��:� ٸ�� �{/�� �{.' ���xz0�(. 	|�zЃb  c3  �X��  :� ~��| H��  AՀ#K��p=� ~=z9� ?}����:� ֈ�: Ј��V b�  :� ֠��P b  : Ш�B ����  
  ~������{.�:�  ��  :�  ��0:` �~P�^����� ��A �� ��! ��1�:���*�� ��� ���$��:~&���bw  :@@@RR�zR �S  �S ;1�و�c8  :�@@R��z� ��  �� :�P9�" =� �����z�' �`�x(2 	|�zw�b�  b�  � :�" >� :@ ?~I��Q�U ":� Ԉ�:�  ר�� b�  :� �p�� b�  :� ט�  "*�F���Io�9i�B ��a�  b�  cb  K�⡂^ʊ>Β^Ϛ>��^�zn��.  -� @�  ;  � ��� ��� ���ʚ��H  :   �> ��Z ��z ��^ʚ~�=� =r:`���(|�b�  b  ���>� ~��;�ꠁ{' �@�x(1 	|�zU�b�  c  �T�AՀ#���| Ha�  ��x�0 ��  Ȉ~��N� >  ���z��:@ �S  ��(=� ~r��{6���  ~7x A�8H  lH  h>  ~��:���@�(|�bX  b�  ��AՀ#K��D>` }ݚ����� ��� �y���0  :� ~Q�|  �~Y4���0  AՀ#K��x?  ~���t��~  ��  -7�A� ��  -�  A� 9����  ��  
  y�  x�:5��z2  ��2�~Y�| H{0d~t��:��.0  z��~�@�   #�3T��r�qS�?:s ט��� b�  K��`n  `�  ).  y� x�| H~� �y�zz1y��{,b#  K��xy `�  >� ~}�:� r�3 p~�*�� �9�" =� 9� p� ��@�y�' � �x(8 	|�z2�bX  a�  � "8� 
a�  ~��b�  N�!ꀁy�' ���x(0 	|�z��b�  a�  ��:@ 
�]  �=  )�  @� |?  }����z����  * @@� `=� ~=z�Q�zp�;0 ـ�� �{4����{5' ���xy��(5 	|�z������  9� ~O�| H�]  AՀ#K����}  )3  A� ��  :� }Ԁ| H>� ~ݪ��{1�~�r׈����z���`�z�' ꀁxzo{(0 	|�z�{a�  b�  ����  )�  @� �?  }����z2��r  * @@� p>� }����z��z��  $]hee^�����};6��; ���� �{.�� �{2' �`�xz0�(2 	|�zp�b  c7  ����  :� �| H�  AՀ#K��p=� ~=r�Q�zy��  � `��  z�  ��9� `a�  c$  b�  K�3�  ~���x��  1� 	| H�� `:Z��r  � � �u  �� `/��x��� `2� | H�� `; ���  ��  :Q�� �zS' ꠁx(3 	|�z��b  bW  ���� `��  �  {  ��bC  a�  a�  K�3�=  ��z��~�И�b  ��  ;  �}��| Hy�  x�:� @b  b�  a�  K�#:� �� �z�' ���x(3 	|�z��c.  b�  ���;  ��  ��  z�  ��b�  bD  b  K�3�  ���z��3�٘�c/  ��  ;  ~��| Hz�  ��:� @c#  b�    %��=0d�ݍ.b  K�#:� ?~���� ���:� �Ԉ�:q ӈ�� b�  :� Ԩ�� bv  :v Ӱ�B ��� �zW' ���x(7 	|�y��b  bY  ��9� ���  ��  )6  A� ��  :� }��| H>@ ~���{1�}�zΈ����y��ꀁy�' ���xz��(5 	|�z��b�  a�  ���]  )�  @� �=� ~=z�Q�zt���  * @@� p>� }ݺ��{6�z��9���: π��@�y���`�y�' ꠁxzr�(4 	|�z��bV  a�  ����  ;  ~�| H�  AՀ#K��p>  ~}�:� ?~�����9� Ϙ�:S Ҙ��� a�  9� �p��� bX  :X ���B ���=  
  0�Ȉ��z��;   �  9�  ��0:� ��P���>��! ��� �� �  &6�*ܳkH(5?���� ����; �~��*�! ��� ���$�>:�&���b�  :�@@Rրz� ��  �� :��՘�b�  ; @@S�{ �  � 9�P:=" >1 ��� �y�' ���x(6 	|�z��c4  a�  �� ;" ? :� ?~������ "9� Θ�;8  ���� a�  9� Έ��� c7  ;7 ٸ�B ��b  c  cb  K��ł�ʊ~Β�Ϛ~����z����  - @�  :� �� �� �� ��ʛ�H  :`  �~ ��� ��� ���ʚ��AՀ#K���`   :   �> H >� ~]�9�P;/ T�x�c.  :�  ��  �� : d�x�b  :`  �p  �p :� y�x�b�  :   �6  :�@���z�' � �x(4 	|�{.sa�  b�  ��r���z��r�: ��*9� 
���:   �2`�2h  '�Z�L�����K�ꀁz�' ���x(9 	|�yԣ���:�  ���:��:`@@Rs�zs ;  	��v  �v 	�v 	B ���v AՀ#K���AՀ#K���A݁�8! � (|�����N� !    ����[�D0        �����������|�� (�!��`[  �A  < D� c�  ;�6@?� ��A݀�B (`|  �;  c>  �>�) A�  ;  �>�;=2?9 c#  cb  H G�H H�>�)� A� H h;  �>�;   �> ?  =�; �>ࣙb���z��f���b��%��  :� ���b�  ; @@S�{ :� ?~���  � 	� 	B ��:� ?~���� ���; ��Ȉ:��Ȉ� c  ; ذ��� b�  :� ט�B ���^�zv�:�  ��  :�  ��0:@ �^P�~���� h�a `�� `�� h��:@�  (�4W���7�J8ܟ~ّ*� `�a h�~$��:�&���b�  :@@@RR�zR �T  �T :y��Ȉbu  :�@@Rրz� ��  �� :^P:�2>� ��ꠁzV' �`�x(6 	|�zu�b�  bQ  � :�2>� :` ?~i���� ":Y�Ȉ:6  Ѱ�� bP  :P Ҁ��� b3  :3 ј�B ��8� b�  cb  K��у>ʊ~Γ>Ϛ~���z����  . @�  ;  �> ��z ��� ��~ʚ��H  :�  �� �� ��� ��ʚ��>� �:8 ��Z ��: ��Q  �1 :q ӈ�bt  :�@@R��z� :  ?~	���  �� 	�� 	B ���� �� :� ?~���� ���
:X ����;8
���� bT  :T Ҡ�� c5  ;5 ٨�B �����z��:�  ��  :�  ��0:  �>P������ x  )�'j�#�P��� p�� p�� x��:`�~��*� p�! x�>$��:�&���b�  :�@@R��z� ��  �� :�����b�  : @@R1�z1 �7  �7 :�P:2> ��ꠁz�' �`�x(6 	|�zu�b�  b�  �� :=2>1 :` ?~i��
�� ":�
���:�  ֈ�� b�  :� ׀��� b�  :� ֘�B ��8� b#  cb  K�ӽ�ʊ~ΓϚ~���z���0  - @�  ;  � ��z ��� ��~ʚ��H  :�  �� �� ��: ��ʚ>Ϋ>(:@ ~ٖ|  �b�  K��`w  `�  b�  c  K��`�  `�  `�  zs  �� �� �}  : 0:0 р�b2  ;  b#  c�  c%  K�3>� ~��� �zT�ꠁzS' � �xz��(3 	|�z�c  bQ  ��;   �= P�� R  *�*�{�
8��r-� @� �>� ~���U�zx��8  * �@� h� R:� ~�����= P>� ~���T�zu�; ب�� �{����{' ���xz�(9 	|�zыb2  c  �T�AՀ#K��x�� V�6) �@� h>� =���z6�z��:v��; ����@�zt�ꠁzw' � �xz��(7 	|�z�bP  bq  ��:� `��  � Dc � D>� ~����� �:] 0� �{6�}���@� $z�' *3 	@� zT' )4 	A� �֐�~��P��:  ~�P|  �
  �  ;  � `;:�:} `��  �Y ��  �S �  :3 ј�2 | H� `z�  ��b#  b�  c  K�3�7 `~��Ԙ��W `2 | H� `:� ��5  �4  :��� �z�' �@�x(9 	|�zX�c  b�  ���� `  +��;7��f�9��  �=  z9  ��b�  bd  c%  K�3�]  ��z��~����b  �}  ;  �~��| Hz�  ��:@ @b  bD  b�  K�#; �� �{' �`�x(9 	|�zq�b4  c  ���:  ��  �]  zY  ��c  b�  c%  K�3�}  ��z5�~��Ԩ�b�  �  ;  ~�| Hz  ��:` @b�  bd  b%  K�#:� ?~��� ��:W �Ҹ�:и�� bS  :S Ҙ��� b  : Ј�B ��� �z�' � �x(8 	|�z9�c4  b�  ���:` ��}  �  )�  A� ��=  :� 6�| H>� ~�����z���ؘ�� �{�� �{' ���xz0�(5 	|�zЃb  c  ����=  *9  @� �>` ~]���z5��  ) @@� p>� ~ݺ��{4�  ,^���g�r-��z��:��:s И��@�z�ꠁz' � �xz��(7 	|�{�bX  b  ���  :` ~3�| H�=  AՀ#K��p>� ~��:  ?~	���:WҸ�:�ָ�� bT  :T Ҡ�� b�  :� ֘�B ���  
  ~������z8�:`  �x  :�  ��0:� ��P��>��! �� ��a �� ��:��~w�*� ��! ��>$��:&���b  :`@@Rs�zs �p  �p :��Ը�b�  :�@@R��z� ��  �� ;P:}2>s ��� �{' ꠁx(1 	|�z��b  c  �� :=2>1 ;  ?	���� ":и�:q  ӈ�� b  : ����� bw  :w Ӹ�B ��c$  b#  cb  K��ق�ʋΒ�ϛ���z���9  -� @�    -³~}4�&�If�:� �� �� ��� ��ʚ��H  :�  �� ��: ��: ��>ʚ>�>� ~]�:r �����Ȓ� �  ; ؘ�c  :�@@R��z� ;  >)���  �� 	�� 	B ���� �� :  ?~)��� ���: �А�:rӐ�� b  : Р�� bu  :u Ө�B �����z��:�  ��  :�  ��0;  �>P������ �� ��� ��� ���: �~�*� ��! ��>$��:�&���b�  :�@@R��z� ��  �� :��א�b�  ; @@S9�{9 �7  �7 :�P;2? ��ꠁz�' � �x(6 	|�z5�b�  b�  �� ;=2?9 :  ?~)���� ":�א�:�  �Ȉ� b�  :� ����� b�  :� ֈ�B ��8� c#  cb  K��ł^ʊ>Β^Ϛ>�  .;S|͙�s�����z���8  . @�  :@ �^ ��: ��� ��>ʚ��H  :�  �� �� ��: ��ʛ>�>` ~�:� ���ЂZؒV ��  :6 Ѱ�b4  :�@@R��z� ;  >	���  �� 	�� 	B ���� �� ;  ?)��P ��P:� �׀�:�ր�� b�  :� ����� b�  :� ֈ�B ����{3�:@  �S  :   �>0:� ��P���� ��� ��! ��A ��P:`�0�*�! ��� ���$�>;&���c  :@@@RR�zR �X  �X ;0�ـ�c3  :�@@R��z� ��  �� :>P:�2>� ���@�z8' �`�x(8 	|�zr�bX  b9  � :�2>� :` ?~i��� ":0р�:U  Ҩ�� b4  :4 Ѡ�� bS  :S Ҙ�B ��8� b�  cb    /^�21�FdvkK�ȱ�ʊ~ΒϚ~���{4���  - @�  :  � ��z �� ��~ʛ�H  ;   �> ��� ��� ���ʚ��>� ~��:W ��: Ԋ ֲ2  � :r Ӑ�bx  ; @@S9�{9 :� ?~���3  �3 	�3 	B ���3 �3 :� ?~��� ��:� �ָ�:WҸ�� b�  :� ֠�� bS  :S Ҙ�B ����z��:   �  :`  �~0;  �>P����� �� �� �� Ȳ: �~��*�a ��! ȳ>$�~:�&���b�  : @@R�z �  � :��ո�b�  ; @@S9�{9 �5  �5 :~P;2? ��� �zt' � �x(4 	|�z0�b  bu  �� ;=2?9 :  ?~)���� ":wӸ�:  �Ȉ� bx  :x ����� b  :   0�@	S�~����Ј�B ��8� c#  cb  K�Ɲ��ʊ>Β�Ϛ>���z���8  -� @�  :� �� ��: ��� ��>ʚ��H  :�  �� �� ��: ��ʛ>�>@ ~ݒ: ��z���� �p  :0 
р�b4  :�@@R��z� ;  >	���  �� 	�� 	B ���� �� �� ;  ?)��V ��V":� �װ�:"а�� b�  :� ����� b  : Ј�B ����{3�:@  �S  :   �>0:� ��P���� ��� ��! ТA زV:`�6�*�! Т� ز�$�>;&���c  :@@@RR�zR �X  �X ;6�ٰ�c3  :�@@R��z� ��  �� :>P:�2>� ���@�z8' �`�x(8 	|�zr�bX  b9  � :�2>� :` ?~i��"� ":6"Ѱ�:U  Ҩ��   1A��t\ClA��eb4  :4 Ѡ�� bS  :S Ҙ�B ��8� 
b�  cb  K�ą��ʊ~Β�Ϛ~���{4���  . @�  :� �� ��z �� ��~ʛ�H  ;   �> ��� ��� ���ʚ���2b  K��`w  b�  K��xr `�  >� ~}�;  r�S p~3�*;3 �:� �Ȉb�  : p��  �� �� ��  �@�z��� �z�' � �x{�(9 	|�z�bV  b�  ���:�  �� P�= R- 	@� �?  =���z���P  )� �@� h�� R:� ~�����} P>  ���z��: �Ȉ�@�z����z' � �xzғ(3 	|�z2�bT  b  ���AՀ#K��x?  ~���� yV�6* �@� h>  ~���z��zX�;2��; ������{6��`�{1' ꀁxzw�(1 	|�z��  2J/��	�%�R߲b�  c5  ���:@ `�Y  � �c �� �>` ~=������ �:� �� �{4�}4��@� $z�' )� 	@� z�' *0 	A� �aԨ�~u�P�a:� ~ӼP|  �
  ��  �  � `�=  {2  Ȉ: `b  b�  bE  K�3�  ~p�Ӏ���  2� | H�� `; ��8  �3  :���@�z�' ���x(5 	|�z�bX  b�  ���� `��  �}  zu  ��b�  b  b�  K�3��  ��{2�~Һ֐�b�  �  :� ��| H{  ��:� @b�  b�  c%  K�#:Q ��`�zU' � �x(5 	|�z�bv  bW  ���;  ��  �=  {5  ȈbC  b�  b�  K�3�  �Q�zw�~ׂָ�b�  �=  :� ~Y�| HzS  ��:  @b�  b  be  K�#:� ?~��� ��&  3�5..Z	O�h��:� �Ո�:Q&҈��� b�  :� Հ��� bS  :S Ҙ�B ��� �z�' �`�x(8 	|�zy�c6  b�  ���:  ��  �  )8  A� ��}  :� 4�| H>� ~ݺ��z8�~X����ꠁzS�ꀁzW' � �xz��(7 	|�z�b�  bQ  ���=  )�  @� �?  ~}����z���T  * @@� p>� ~=���{0�z�:p��:� Ӱ����zt��@�zu' � �xzW�(5 	|�{�b�  by  ���  :� ~��| H��  AՀ#K��p>@ ~��:` ?~i���&��*;5&٨�;*ب�� c4  ;4 ٠�� c  ; ؐ�B ���}  
  ~w�����z6�:@  �V  :�  ��0:` �~P��>��! �� ��A �� ���:��~U�*�a �! �  4vV����M`c��>$�~:&���b  :@@@RR�zR �P  �P :��Ԩ�b�  :`@@Rs�zs �t  �t :�P:]2>R ��� �z�' �`�x(1 	|�zp�b  b�  �� :�2>� :  ?~)��U*�T ":�*֨�:  Р��� b�  :� ֈ��� b  : И�B ��b�  b�  cb  K��݂^ʊ�Β^Ϛ���^�zq���  - @�  9� �� ��� ��� ���ʚ��H  :�  �� ��Z ��z ��^ʚ~�>  }��; ��:���8  � :� ���b�  :�@@R��z� :� ?~����  �� 	�� 	B ���� :� ?~���O ��O.:/ ��x�;/.�x��� b0  :0 р��� c8  ;8 ���B ����z��:`  �n  :@  �^0;  �P������� �� ����  5(�W��1Pu�:��~ϩ*�a ����$�~:^&���bX  :�@@R��z� ��  �� :��x�b  :�@@Rրz� ��  �� :�P9�2=� ���`�z�' ���x(8 	|�z�bv  b�  �� :]2>R :� ?~���.�� ":.�x�;  ؐ��� b  : И��� c  ; �p�B ��8� bC  cb  K��͂�ʊ�Β�Ϛ�����y����  -� @�  :� �� ��Z ��� ��^ʚ��H  :�  �� ��� ��� ���ʙ��:`  �~ H <>� =�:9`; T؈�c  :�  ��  �� :Q d҈�bU  :�  ��  �� 9� yΈ�a�  :`  �n  :�@� �z�' � �x(6 	|�{�b  b�  ����Z��: �9�9��~Yy*�z������y�:��� �z�' ꠁx(0 	|�  6������v��c3z��c  b�  �b:� ���:@  �Yp�Yx���z�' �`�x(. 	|�zo{a�  b�  ���:��; @@S�{ :  ~)��  � 	� 	B ��� AՀ#K��AՀ#K��A݁�8!`� (|�����N� !        ����[�D�����!���A��|�� (�!�A`[  �A  < D� c�  ;��?� ��A݀�B (`|  �;  c>  �>�) A�  ;  �>�;=�?9 c#  cb  H )aH 4�>�)� A� H T;  �>�;   �> �> �8�Ȉ���z��:�  ��  :�  ��0:� ��P�>`��h�� h�! `>� ~���! `�� h���:��7�*�! `�� h��$�>:�&���b�  ; @@S9�{9 �6  �6 ;7�ٸ�c6  :�@@R��z� ��  �� :�P:��>� ��  70q�7N�PD � �z�' ꀁx(5 	|�z��c4  b�  �� �� H;=�?9 � @c  c#  ~��b�  N�!`t  b�  �� ��ʋ>Γϛ>���z���  . @�  ;  �> ��� ��� ���ʚ��H  :�  �� �� ��� ��ʚ���� �-7��;  A� ;   -�  A����z��;   �  :�  ��0;   �>P�0��8�� x�� p?  ~���� p�! x�6�:��~��*� p� x�$��;>&���c7  :�@@R��z� ��  �� ;�ذ�c  :�@@R��z� ��  �� :�P;=�?9 ��ꀁz�' � �x(7 	|�{��� :��>� ; ꠁ{�� �{' �`�x{5�(4 	|�zu�b�  c  �W b�  cb  H �;  )�� �� ":v  Ӱ��� c  ; ؐ�  8�\l.��`�מ�� by  :y �ȈB ����ʊ�Β�Ϛ�����z���Y  . @�  :� �� ��� ��� ���ʚ��H  :�  �� ��: ��Z ��>ʚ^�:z ��xs A� �  �� ��  �� H  �� �� ;= ��c2  ?  ~��:�  :` �c#  b�  be  K�3:� ~��c�  :U �Ҩ��  �  � 	� 	B ���:(��,�z.�5  �� �u :� ר�b�  ; @@S��  � :� ��:�� �� �6  :v 
Ӱ�br  ; @@S�{ �  � :� :� @��  ;7 ٸ�c2  ; @@�  S�� �^�zt�;   �  ;   �>0:@ �^P�~ �� ��a �� ��! ��5�:@�~��*� ��a ��~$�;>&���c4  :@@@RR�zR �Y  �Y :u�Ө�bx  :�@@  9/������R��z� ��  �� :^P;=�?9 ��� �zT' �`�x(4 	|�zx�c  bQ  � :��>� :u ��@�z�' � �x(8 	|�z2�bX  b�  � "� �z�' ꠁx(1 	|�z��b  b�  � 2�@�z�' ꠁx(1 	|�z��bX  b�  � B���zp' � �x(0 	|�z6�b�  by  � Rb�  cb  H I��ʊ�Β�Ϛ����z2��r  - @�  :� �� ��: �� ��>ʛ�H  :�  �� ��� ��� ���ʚ��:   � :   �> H <>@ ~}�:�P;6 Tٰ�c8  :�  ��  �� :� dհ�b�  :   �  � :6 yѰ�b2  ;   �  :�@� �z�' � �x(7 	|�z�c0  b�  �r�(��0���:@�~��*�8��@�� �� �;3 �� �{0'   :�Cy��$@Z!�1���x(0 	|�zыb6  c7  ��R:� ���:@  �S`�Sh� �z�' � �x(0 	|�{8�c  b�  ��:� �:�@@Rրz� :� ~����  �� 	�� 	B ���� AՀ#K���AՀ#K���A݁�8!�� (|����N� !    ����[�D�        �����������|�� (�!��`\  �A  < D� 3��| �A݀�b (`}  �\  c^  �^�) A� ;@ �^�;_��cC  c�  H !]H 
��^�)� A� H $;@ �^�;@  �^ ;@x�_��;_��? ��c9��{9�g9��c9���:  ;: �Јc:  ;@@@�Y  ;_�@;  \�:  ;: �Јc:  ;@@@SZ�{Z �Y  �Y �Y �Y ;_�`;  @�:  ;: �Јc:  ;@@@SZ�{Z �Y  �Y �Y �Y ��{:�;   �  ;     ;�߅
��F+-���>0�У^س^$��>�^��^.; &>�*�^�>$�?�"; �_�*; &>�*�^.�_��?��/x:�x�N   @� \;>����;R����Y  �� �� �� �9 �� �8 �X  �� �� :� ;>Pb�  c$  蠁0���09@ %D A��/�� �;^�� �{U' � �x(5 	|�{8�c  cW  ����:��`� �z�' � �x(: 	|�{�c6  b�  ����;_�@� �{U' � �x(5 	|�{8�c  cW  ����:���� �z�' � �x(: 	|�{�c6  b�  ����;_��� �|�c  cU  ���;?�0���{6' �@�x(6 	|�{W�b�  c5  ���; `��:��;_� ;?��:���:���:����� �X �8 ��  �� (�� 0:� ��  �� c  8� �8�  D  �^ʋ>�  <���2�|k��͓^ϛ>����z����  - @�  ;  � ��[ ��; ��^ʛ>�H  :�  �� ��� ��� ���ʚ��:�H� �(|�c  b�  ���r;_��� �{U' ꀁx(5 	|�z��c6  cW  ����AՀ#��r| Hb�  �[`�8 ��  Ȉ~��N� ���z��;   �  ���{:���  )� �A�`H  XH  T:�hꠁ(|�b�  b�  ��rAՀ#K��h������ �� �z���:  3 | H{ ����  AՀ#K�������2� | H
  �������b�  �! �?�����.8 A� ����-7 @� L�\ �:���:���� �� �z�' ���x(9 	|�z��c  b�  �V "8� db�  ~��cB  N�!;  �� ~��P|  �b�  �:` ~X�|  ��_������-� A� ���.5  @� L�\ �;?��  =KG�v/�jl�:���� ��`�z�' ���x(2 	|�zӛbp  b�  � "8� dc#  ~��cB  N�!�:� ����:_��-8  zV�~��@� :� װ�b�  �a� �zp�� �zt' �@�x{1�(4 	|�{Q�b4  bu  �������)� @� �_���_��H  :� �����a�����������z  ��;_��bc  cD  c%  K�3�?�����z��~X����bV  �������~w�| Hzz  ��;  @bC  c$  cE  K�#AՀ#K������b�  K��xu �b�  K�|q���?��;   ���:� ����: 3�� :�  ���:`  �� :@ �_�0��{:�:�  ��  :�  ��0�>P��X��$�>�p��x��.:`&~�*�^�$��"; �~_�*:�&~��*�^.�_�����x6�x�  >fs�7�5,ժ��iN   @� \:>P���:�R����  �q � �Q �1 �W �7 �  �w � ;^ :�PcC  b�  蠁0���09@ %D A�� �:������z�' � �x(2 	|�{6�b�  b�  �_��;�����{' ꠁx(: 	|�z��b�  c  ���;?��ꀁ{6' �`�x(6 	|�zt�b�  c7  ����:_���@�zU' � �x(5 	|�{�cP  bQ  ���:�0� �zt' ���x(4 	|�z��c4  bu  ���:�� � �z�' �@�x(2 	|�{X�c  b�  ��:���`�z�' ꠁx(9 	|�z��bp  b�  ��":�� �@�z�' ���x(: 	|�zғbX  b�  ��2:������z�' � �x(3 	|�z7�b�  b�  ��B:���@�z' ꀁx(6 	|�z��cR  b  �_�R:?��ꠁ  ?�K�]�|���1�z7' � �x(7 	|�{5�b�  b3  �_�b;�����|�b�  c  ��r:� `��;_�p:��`;?�P:��@:�0:_� ;�:�� :?��:��9���9����T �� �4 ��  �t (�T 0� 8�� @�4 H� P�� X�� `;@ �T  �T b�  8� �8�  D  ��ʋ>Β�ϛ>���z���S  - @�  ;  � ��� ��; ���ʚ>�H  :   � ��� ��� ���ʙ��;] ���� z��:� ~��:����u  �y  �u 	�y 	B ��:@ �_��H  ;   � �?��)� A� L� �9���9����� ��@�y�' ꀁx(7 	|�z��cX  a�  � "8� �a�  ~��b  N�!H �:`  ���:���:U TҨ�bQ  :�  ��  �� :� dԨ�b�  ;@  �T  �T ;5 y٨�c8  9�  ��    @Th�m&���K�x�:�@� �z�' � �x(3 	|�z0�b  b�  ��������[��_��9���~�q*�[��������������_��;?���`�{1' � �x(1 	|�z�bt  c5  ����:@ �_��:�  �����������z�' ���x(8 	|�y�sa�  b�  ��;_�0; @@S9�{9 :` ~i��:  �: 	�: 	B ��:���:���:@ ~I���  �� 	�� 	B ���� :���; ��9� }���  � 	� 	B ��� :�  ����9�  ����:?��: @@R�z �  � :` @���AՀ#K���AՀ#K���A݁�8!`� (|�����N� !        ����[�D�����!���A��|�� (�!�A`[  �A  < D� c�  ;� ?� ��A݀�B (`|  �;  c>  �>�) A�  ;  �>�;=�?9 c#  cb    A�q>�r�C��=2H �H �>�)� A� H �;  �>�;   �> ��{8�;   �8  ;   �>0���>��! h� `?  ��! `�� h���:��8�*�! `�� h��$�>:�&���b�  ; @@S9�{9 �7  �7 ;8����c7  ; @@S�{ �  � �� �;�? �; �c  )�b�  N�!;�? ��;8 ����� z��� ���ʋ>Β�ϛ>����z����  . @�  :� �� ��: ��� ��>ʚ��H  ;   � ��� ��: ���ʛ>�>� �����! �{6����{5' ꀁxz׻(5 	|�z��b�  c5  ����z��� b�  K��`t  �� z���� :� ;:�c�  8� 
b�  8� 
c'  9  K��ꠁ|�b�  c�  �� b:� 
��  �=  )9  @� �  B��D�V|&�L>� ~��� f{6���  )� @@� h>� ��� fz��:� �Ȉꠁz�����z�' ���xz��(9 	|�zիb�  b�  �� b�=  :� ~��| H��  AՀ#K��x��  *7  A� ���  ;  8�| H>� ~���� fz��~��������z��� �z�' ���x{6�(8 	|�z��b�  b�  � r��  )7  @� �>� ~ݢ� v{5���  )� @@� p>� �� vz��z��:���;9 �Ȉꀁz�����z�' ꠁxzԣ(9 	|�z��b�  b�  �X r��  ;  ~��| H��  AՀ#K��p>� ~���T fzx���  �� 0�=  {5  Ȉ:� 0b�  c  b�  K�3�]  ~w�Ӹ���  36 | H�4 0;���  �X ��  �S ��z��� ����^�zv�:�    C�����������  ;   �>0;  �P�^��~��a x�A p�� p�� x���; �~��*� p�a x�~$�:^&���bV  :�@@R��z� ��  �� ;4�٠�c3  ; @@S�{ �  � :�P:��>� ���@�z�' �`�x(4 	|�zr�bX  b�  � �:}�>s �� b�  bc  ~��b�  N�!:W Ҹ�� {5��� ��~ʊ�Β~Ϛ�����z���  . @�  :@ �^ ��: ��z ��>ʚ~�H  :�  �� ��� ��� ���ʚ��� �;   �  >@ =��`�z�����z�' � �xz�(4 	|�{�bv  b�  �� b�]  )2��@� D�  ?  ~���U fzw�~עָ��6  )�  A� �  2X | H�]  AՀ#K���>� ~}�� 0:� 0~עָ�b�  �! �� f  D��� �)ջ����z��� ��S 0:���z� ~Ҹ| H�  �� @�� P� P�� @~7�@A� >@ ~���� P�� @>` ~���� @�! �� ��U 0~Ҹ| H�� 0z�  ��c#  c  b�  K�3:u ��@�zv' ���x(6 	|�z��U b�5 0)9 �@� ?  ~��:� ��� @H  >� ~}��S 0�S @>� =�� @�  ��  z�  ��:� 0:Y �bC  b�  b�  K�3�}  � fz��~ؚ���b�  ��  :� �~��| Hz�  ��;  @b�  c  be  K�#:\ ����� z��:� ~���Y ��T ; ��Ȉ�� c  ; ب��� b�  :� Ԙ�B ��:@ �Y H  :`  �~ >� ~���� )� A� X�[ �;=�?9 >� �:x � ����zv' ꀁx(6 	|�z��b�  bq  � "  E�'� S�e �R8� �c#  ~��bB  N�!H  �?  ~��:�  �� :v :� Tט�b�  :   �  � ;3 d٘�c5  :@  �Y  �Y ; yؘ�c  :   �8  :@���z' �@�x(5 	|�zW�b�  b  �B�z�������: �~v�*:� 
��p:@  �V0�V8���z' � �x(9 	|�{�b�  b  �V�:�  ����AՀ#K��AՀ#K��A݁�8!�� (|����N� !    ����[�D�        ����!���A��|�� (�!��`[  �A  < D� c�  ;�@?� ��A݀�B (`|  �;  c>  �>�) A�  ;  �>�;=?9 c#  cb  H 
�H 	��>�)� A� H 
�;  �>�;   �> � O� �?  ��� ��� �;: �� �z����  ��  ~6�@;   A�   F�'p'Y;�; ��A� ;  � �= -  A� :� ��  H  L:� ?  =�� �z��� ��  �7 �� }��@@� }��@A� :� ��  H  :�  ��  �  .4  A� �?  ~��;5@���{6' ꀁx(6 	|�z��b�  c3  �U ��� Fz��:� ��  �}  zr  ��c#  c  bE  K�3:�����z�' �`�x(4 	|�zw�b�  b�  � ��\ Vzt�:� ���  �=  {8  Ȉb�  b�  c  K�3H :�  �� �\ /�A �>� =�� ��� �:�(�A �zx���  ��  �� �6 }7�@@� �� �� }4�@@� }7�@:@  A� :@��A� :@ �] �} -�  A� ;   �  H  L:� ?  ~���T �zu��� �  �5 	�V ~7�@@� ~9�@@� :� ��  H  :`  �}    GE�k��e�k�;�  -5  A��>� �����Zċ:ƒ�@�XD�8F�\ ?�X �:� ��  �  )�  A� ���  :� 7�| H>` ~]�� �z��~��������z��ꀁz�' � �xz��(5 	|�{7�b�  b�  �� ��  *8  @� �>` =��� �z����  ) @@� p>@ ��X �zv�z��:���;9 �Ȉꠁz���@�z�' ���xzU�(3 	|�zիb�  b�  �X ��=  :� ~��| H��  AՀ#K��p>� ~���U �zx�;  �5 0:��:� 0��  �T ��  �V �}  ;6 ٰ�2� | H�� 0zw  ��c#  c  b�  K�3�U 0~��԰��u 033 | H�5 0;���  �X ��  �T �u 06�ٰ��� Vz���U 02� �| H�� 0:` �c#  c  be  K�3:��  H�E�Y G�g;<����z�' ꀁx(2 	|�z��b�  b�  � ��u 0)� �@� >@ ~��:� ��� @H  >� =�� 0� @>� ~}��S @�]  ��  z�  ��:� 0;�c  b�  b�  K�3�=  � �z��~��֐�b�  ��  :� �~w�| Hzu  ��;  @b�  c$  b�  K�#H  h:@  �^ ?  ~��:���`�z�' � �x(6 	|�{3�bx  b�  � �� Vz��:� ���  �}  zy  ��b�  bD  c%  K�3;   � :�  �� >� ~ݪ:v ���ЂZأ:ܒS �3 ��  ; ؘ�c  :�@@��  R���� :@ ��V P� &{7��� �:v ���ࢺ�Z撓  �� �S ; ؘ�c  :�@@R��z� :� ~����  �� 	�� 	B ���� :@ �V `:v p;  @�3  :�   I2w��߶7�^�;�՘�b�  ; @@S��  � ��{2�:`  �r  :�  ��0�����$���>��~��~.:@&>�*��$�:��~��*:`&~~�*�>.�6��v��x2�x�N   @� \;����;>R����x  �� � �� �X �� �Y �y  �� �� :�;Pb�  c  蠁0���09@ %D A�^�A ��� �:��>� ~��� �z�' �`�x(8 	|�zy�c2  b�  �UR:� p� �z�' � �x(4 	|�{8�c  b�  �Ub:� `� �z�' � �x(6 	|�{�c2  b�  �Ur:� �� �z�' � �x(4 	|�{8�c  b�  �U�ꀁz�����z�' �`�xzԣ(8 	|�zt�b�  b�  ��:U P���zS' ���x(3 	|�z��b�  bY  ��:���`�z�'   JTaٮ�������@�x(7 	|�zS�bx  b�  ��:� ����z�' ꀁx(2 	|�z��b�  b�  �U�;5@� �{4' ���x(4 	|�z����:� `��:u�:U�:��:��;5�;�:5p:`:�P�w �W �� ��  �7 (� 0�7 8� @�� H:` 	�w  �w b�  8� �8�  D  �^ʊ�Β^Ϛ����{6��6  - @�  :  � ��� ��z ���ʚ~�H  :�  �� ��Z ��� ��^ʚ��;   � H ?  ~��:6`: TЈ�b  :`  �p  �p :� d׈�b�  :�  ��  �� ; y؈�c  :�  ��  :~@� �zr' ꀁx(2 	|�z��b  by  �����:�6�:��~��*:@ 
�V�:�  ��p��x� �zy' � �x(9 	|�{�b  bu  ���:6@:�@@  K�A������0�aɲ�  R���� �� :V�; @@S9�{9 ;  	��2  �2 	�2 	B ���2 AՀ#K��hAՀ#K��pA݁�8! � (|����N� !        ����[�D@        �A���a�����|�� (�!��`\  �A  < D� 3� | �A݀�b (`}  �\  c^  �^��^ (;@  �^�;@  �^�^ *-  A��^ *-� A���^ *. @� ;@ �^H  �^ *- @� �;@ �^�^  �A H  �;^P;;�� �(|�� H �;>�;��@�(|�cV  c  �� H �;P;[����(|�b�  cU  �� AՀ#��| Hc6  �[�� �  ��~��N� H  4�A )�  AՀ#A����A * AՀ#A��d�A ) AՀ#A���:�  ��H !��> *-� A�!H�
.  A� \  L��armxLN
}���z��;@ �U  �;?�`;@�����{' ꠁx(: 	|�z��b�  c  �Y "8�"�c#  ~��b�  N�!;@ �^�:�� �(|�c  b�  ��RH ��] /�^�� ?��� O����� _����] o�^r� �b� ���R�� ���B�] ��^2� ��"� ����� ����] ��^�� ������ҋ^) @� l:�  ���:�0�`�(|�bx  b�  �bH �\(:��`:�@�\ ���z�' �`�x(6 	|�zw�b�  b�  � "b�  I�bB  N�!��)�  @� ��] zt��� b�  K��xy �� �`{5�"S5&6S5.S5#~��xz� ���z���^���tH  $:������t�[܊{�zSB,�~�zt�����?�vc#  K��xx �ꠁ`{�"S&6  M�����H�Q`S�S.S#Z�x{Z �^�{W����:� ���^* @� �:~)`ꀁzy' � �x(9 	|�{�b�  bw  ���:���@�z�' � �x(2 	|�{:�cR  b�  �^)�� �z�' ���x(4 	|�z��c  b�  �^)�:� ��9;  �>+C;[Hꀁ(|�b�  cW  ��*:� ����) @� :`  �~:@  �^H �;>�;Y ��ȈcT  :�@@R��z� ��  �� �� �� ��  �� ":� ��Ȉb�  ; @@S��  :y �Ȉbr  :���R����  �� ��)� @� ;@  �^H  H  � *.  A� ? \�c��{�g�@c@@��>�\�b���z��f���b�@@���;   �> �:@ �^����) �@� (:~����bw  ;@��SZ�{Z �S  �S H @:�����b�    N��y�N��:�.:���Rրz� ��  �� �>�)� �@� :@  �^�H x:� �� e* A��^�) �A��:` �~ eH ���-�aA� ����.fA� ���z���� �x2�x�M   A� T�^�zz�� �z��:�`���(|��� ��{2�AՀ#� �| Hb�  �[�� ��  ��~��N� AՀ#�| Hc5  ��U �u  ��~i�N� ����� ���{:�� ����^�zv�� �x7�x�M�  A� ,��z���Z �zy�;x���(|�b�  c  �� :��`b�  c�  H UAՀ#�^| Hbz  ��� �  ��~��N� ���� ��<8:��`:~@�\0�@�zv' � �x(6 	|�{�cT  bu  �� ":�  �� 0�� 8b�  ~I�c"  N�!H  ? \�c��{�  O\-1l�����g�@c@@�܊~�* �A��?@\�cZ��{Z�gZ@@cZ@@�^�H �:�*�~��*���}4�@@� ��+�[�}7�@@� �;;��  �Y{ "�~U;^ ꠁ{V' ꀁx(6 	|�z��b�  cW  ��)�:[�� �(|�c4  bU  ��)�;   �+6H L�^)�zz��� ��r�v{5���  :^ ���  �^vzz�:� �Ј:�	 ;  	��7  �6  �7 	�6 	B ���� �� �� �� AՀ#�^R| Hbz  ��: ��  Ȉ~��N� ��������:��>:��� �:`�~��^�-� d@� p�^0�^��>*�*��v:�n>�*:�::��:�:���:~�����V  �S  �V �S �V �S �V �S �V  � "�S  � "�>|�>#����� �:�  ����:��`b�  c�  H �  P����)�D_AՀ#�^R| Hbv  �[� �6  ��)�N� >�\�b���z��f��@b�@@�����z��:@  �S  :�  ��0;   �P�^��>ȳ! h�A `�� `�� h���:��~��*�A `�a h�~$�^:�&���b�  ; @@S9�{9 �6  �6 ;^����cT  :�@@R��z� ��  �� :�P:��:S�Ҙ�� �z�' ���x(9 	|�z��c  b�  �� :��`b�  c�  K�a̓^ʊ~Γ^Ϛ~���{5���  . @�  :� �� ��[ ��� ��^ʚ��H  ;@  �^ ��{ �� ��~ʛ��v{5�:� ~��:����U  �V  �U 	�V 	B ���� �� �^�zz�;   �  ;   �>0:� ��P����� x�� p�� p�A x�^�:`�~ޙ*� p�A x�^$�;>&���c7    Qi~j-�)�zl$d:�@@R��z� ��  �� :�����b�  :�@@Rրz� ��  �� :~P;_��;��Ј���zt' � �x(4 	|�{7�b�  bu  �� :_�`:� ~��;_��;2  ِ��z  �y  �z 	�y 	B ���� �� bC  c�  K�j]��ʊ�Β�Ϛ���^�zx���  - @�  ;@ �^ ��� ��; ���ʛ>�H  :�  �� ��� ��[ ���ʚ^��^�zx�:�  ��  ;@  �^0:�  ��P�>P��X�� ��! �� ��A ��^�:`�~��*�� �� ��$��;^&���cW  :�@@R��z� ��  �� ;>����c2  :�@@R��z� ��  �� :~P;��:��������zu' �@�x(5 	|�{W�b�  by  � :_�`:���ꠁz���`�z�' � �xzu�(7 	|�{5�b�  b�  ��   R7B�h^g�YC0nbC  c�  K�й;  	��T �_�;_� � b�  :� Ԩ�� cW  ;W ڸ�B ����ʊ~Β�Ϛ~����z����  -� @�  ;  �> �� ��{ ��ʚ~�H  :�  �� ��� ��[ ���ʚ^�:�
0�@�z�' � �x(4 	|�{:�cR  b�  �_�;  �������z�  ��:�� b�  b�  b�  K�3��{:�:��Z  �� �� �S  :� 
՘�b�  :�@@R��z� ;  	���  �� 	�� 	B ���� ������_�/bX  by  �����?b�  b�  ����Ob�  b�  ��"�_�_bX  by  ��2���ob�  b�  ��B�_�p�_�P��z��:@  �S  :�  ��0:� ��P�>@�H� ��! ��A ��� ����:��^�*�A ��a ��~$�^:�&���b�  ; @@  S��!�˻��D�-S�{ �  � ;>����c4  ;@@@SZ�{Z �Y  �Y :�P:��:S�Ҙ����z�' ���x(8 	|�z��b�  b�  � :��`�_���T "���b�  b�  �T 2��c  c3  �T B���/b�  b�  �T R��?c  c3  �T b���Ob�  b�  �T r�_�P�T �b�  c�  K��1��ʋ>Β�ϛ>����z���x  . @�  :@ �^ ��[ ��� ��^ʚ��H  :�  �� ��; ��� ��>ʚ�����z��:`  �x  :@  �^0;@  �^P� ��(�� ��� ��! ��� ����:��>�*�a �� ��$�~:^&���bZ  :�@@R��z� ��  �� :�����b�  ; @@S9�{9 �4  �4 :�P;��:x�����@�z�' �@�x(5 	|�zZ�cX  b�  � :��`b�  c�    T�$�a�4����'K�ց��ʊ�Β�Ϛ�����z���R  - @�  ;  �> �� ��{ ��ʚ~�H  :�  �� ��� ��� ���ʚ�����z��;@  �R  ;   �>0;   �P�~������ ��a �� ��� ����:��~��*�A ��A ��^$�^;>&���c8  :�@@R��z� ��  �� :~����bv  :�@@R��z� ��  �� :�P:_��;R�ڐ�� �z�' � �x(4 	|�{8�c  b�  �� :��`b�  c�  K�aт~ʊ^Β~Ϛ^���{7���  -� @�  :� �� ��[ ��� ��^ʚ��H  :`  �~ ��[ �� ��^ʛ���{7�:�  ��  :�  ��0;@  �^P��Т~زa ��� ��A �� ȳ�; �~^�*� ��� Ȳ�$��:�&���b�  :`@@Rs�zs �t  �t   U�?�妕"��r��:�����b�  :@@@RR�zR �V  �V ;>P:���:��ո��@�{3' ꀁx(3 	|�z��cV  c7  �� ;�`c  c�  K��Q�^ʊ~Β^Ϛ~���{4��T  . @�  :� �� ��� ��� ���ʚ��H  :@  �^ ��{ �� ��~ʛ���{4�;@  �T  :�  ��0:�  ��P�`�^h�A ��� ��a У س�; �~~�*�A Т� ز�$�^:�&���b�  :@@@RR�zR �W  �W :�����b�  :`@@Rs�zs �u  �u ;>P:���;T�ڠ����{2' ���x(2 	|�z��b�  c3  �Z ;�`c  c�  K����ʊ�Β�Ϛ�����z���y  - @�  :@ �^ ��[ �� ��^ʛ�H  :�  �� ��� ��� ���ʚ�����z��:`  �y  :@    Vk����v���q��^0;@  �^P�p��x�� �� �� �� ���:��~��*�a �! �>$�~:^&���bZ  :�@@R��z� ��  �� ;����c  :�@@R��z� ��  �� :�P;?��:y��Ȉ�@�z�' �@�x(5 	|�zZ�cX  b�  � :��`b�  c�  K���ʊ�Β�Ϛ�����z���R  -� @�  ;  �> �� ��{ ��ʚ~�H  :�  �� ��� ��� ���ʚ��:� ���H |AՀ#K��X>@\�bR��zR�fR�@bR@@�^�AՀ#K��^+C* �@� ��;��ē>:�>:` �~ �:� �����- d@� p��0�����*�^*��^v;@n~��*; :; �:~:���:������  ��  � �� � �� � �� ��  �S "��  �T "��|��#H L�^+�>  W���ˍgC����+�� }��@@� }��@A� $�^�zv�� 0�� 8��+��+���)���z���Z . @� ��^��A ��� �z��� � z��-8  {S�~Z�@� :s Ҙ����zW�ꀁzU' � �xz��(5 	|�{�b�  bU  �� �Y :` ~��P|  �~�4��� :@ �^+4H  lH  h��H:��`:�@:~ ��\@���z�' � �x(8 	|�{7�b�  b�  � "�@�zt' ���x(4 	|�z��U 2b�  I�b�  N�!AՀ#��| Hc4  ���t �T  ��~I�N� :��`b�  c�  H 
MAՀ#�| Hc:  ��� �z  ��~i�N� ���)� �@� H  H  H  H:@ �^�H  <:��� �(|�c2  b�  �^�H 0;��@�(|�cV  c  ���H ���  X펁�l'�?u��f. @� ���- @� \�> �-� �@� P�|:_�`;@�\���{' ꀁx(6 	|�z��b�  c  �� "8� �bC  I�bb  N�!H  L�<:��`;@��ꠁ{' �@�x(4 	|�zU�b�  c  �V "8�#)b�  ~��c"  N�!H  T;@  �^���* �@� ;  ��:� ��H  :`  �~�:@  �^���~�4����{:���  H �AՀ#��| Hb�  �[�� �  ��	�N� ;  �> :�0�@�z�' ꀁx(5 	|�z��cR  b�  �^)b:�  ��)p��)x;�� �{' ꀁx(5 	|�z��c6  c  ��)�;@  �^)��^)�:`  �~)��~)�:@  �^)��^)�:�  ��)���)�:�  ��)���)�;   �)��)�;   �>* �>*:�  ��*��*:�  ��*   Y�/J���dr
�J��*(;@  �^*0�^*8:`  �~*P�~*X:@  �^*@�^*H:�  ��*`��*h:�  ��*p��*x;   �*��*�;  )�:���؈:�*�����W  �V  �W 	�V 	B ��:`  �~+`�~+h:^�ꠁzT' � �x(4 	|�{�b�  bY  ��:�  �� q;@ 1I�:���؈:~�����  ��  � 	�� 	B ��:^�:��Ր�b�  ; @@S�{ �  � � � � :�  �� d;@  �^ e:`  �~ h:� � p:� �� r:@  �^ �;   �>1;   �2:��:� \֨�b�  :`@@Rs�zs �v  �v :� fԨ�b�  :@@@RR�zR �T  �T ;;
� �(|���;[
0�`�(|�bt  cU  ��2:�
H���(|�b�  b�  �B:@  �^��^�;@  �^�:`  �~�:� :���R��z�   Z�̔�K]� ���:� 
~����  �� 	�� 	B ���� �� �� :� ���;  	)�;
`�؈:^0����X  �R  �X 	�R 	B ���{H�~ �:�  �� �:� @�� �:�  �� �:��; @@S9�{9 �7  �7 �7 :@  �^ ;^	 ; @@S�{ :` ~i��  � 	� 	B ��� � � :�����b�  8��K�S>� ���:� ��;  @�>:� ��:@  �^:`  �~;%p���c  8��K�S;@  �^:�  ��:�	�:�@@R��z� ;  )���  �� 	�� 	B ���� :��:@@@RR�zR �W  �W :` �~; �� ;^
0:�@@Rրz� ;  )���  �� 	�� 	B ���� :�  ��$��H�[Lz���^ mzW��� i:`  �~&;  �(;   �>,:�  ��0;@  �^   [@��m��?�8��^:�  ����:�  �� ��(:@  �^0�^8AՀ#��b| Hb�  ��3 �S  ȈI�N� AՀ#�R| Hb�  ���� �r  ��~i�N� ; 
�; :;[
��؈:�:����  ��  � �� � �� � �� �Z  �� "�U  �� "��+?) �@� :~)`� �zx' ꀁx(8 	|�z��c4  bu  ���;@  �^�:@ �^ �� �:��`;@�| �� �{' ꀁx(5 	|�z��c4  c  �� "8� �b�  ~i�b�  N�!;^��@�{X' � �x(8 	|�{2�bT  cU  ��)����{S' ���x(3 	|�z׻b�  cY  �)��^�-� dA� (���� �:�  ����:�`bc  c�  H �AՀ#���| Hb�  �;� �Z  ��~I�N� :�
�:�::{
��؈  \qX@f��DzZ��:�:�����  ��  �� �� �� �� �� �� �S  � "�W  � "�>+?* �@� �:^)`ꠁzT' ���x(4 	|�zիb�  bW  ���:`  �~�;@ �^ � �;?�`:�@�\ �ꠁz�' ���x(7 	|�zիb�  b�  �� "8� �c#  ~I�c  N�!:~��@�zt' ꠁx(4 	|�z��cV  bw  ��)�� �zr' � �x(2 	|�{�c4  bu  ��)�AՀ#���| Hb�  �[� �z  ��~i�N� ;  �>:�
�ꀁ(|����AՀ#K������- @� �^�zv�;@ �V  H  ��{5�:� ��  H  �� ��� �A݁�8!@� (|��A��N� !        ����[�Dx��� ������|�� (�!��`\  �A  < D� 3� @| �A݀`}  �|  c~    ]H���m�K�o��|;_��;>@� ������{5' ꀁx(5 	|�z��b�  c5  �� "c  cC  ~��cb  N�!A݁�8!`� (|���N� !        ����[�D!�      [�D "�       T   H �       	�    [�D1                   (        , �  `#     �6    �#     <     P     |     �     �     �     �          4     x#     �#     �     �     �                D     X     �     �     	     	     	<6    	T6    	l6         [�D -        T   H �        �    [�D1�                ^bFϢ��N?��8     (      O  4     �7    6    \     �     �6    6    T     �     �6    �     4     `6    t     |     �7    7    47         D     �7    �7    �7    7    <7    d7    �7    �7    7    �6    �6    	P7    	p7    	�7    
x#     7    $7    L7    �7    �7    �7    p6    �6    \6    (6    X6    �6    �7    7    <7    �     �     �     �     �     �     �     7    87    `7    P     �7     _�p~��_��b�� �7    7    �7    �7    �7    L6    �6    06    �6    ,6    X6    �7    �7    7    \6    t6    �6         [�D F�       T   H �       (    [�D20                   (        4     �      �     7    $7    H7    �     �     @7    `7    �7    �7    t     7    $7    L7    �7    �7    x6    �6    �     �     �     �     6    ,6    D6         [�D N        T   H �        PP    [�D2�                `�u�S�B�`k��     (     �  4     �6    7    7     7    07    �7    �7    �7    7    $7    47    D7    �6    7     7    07    @7    �7    �7    �7    ,7    47    D7    T7    �     �     6    D7    L7    \7    l7    �7    �7    7    X7    `7    p7    �7    6    X7    `7    p7    �7    �7     7    (7    l7    t7    �7    �7    �6    (6    P6    h6    �6    �6    7    7    $7    47    �7     a�*K�X1��� �7    �7     7    (7    87    H7    �6    6    `7    h7    x7    �7    �7    7    07    t7    |7    �7    �7    7    �6    �           6    �6    �      6    (     4     P6    \     x6    �     �     �6              `     �6    �     �     �7    �7    �7    �7    H     X6    �6         D7    L7    \7    l7    x     �     �7    �7    $7    h7    p7    �7    �7     6    h7     b(w�`&\���g� p7    �7    �7    �7    7    87    |7    �7    �7    �7    <6    �7    �7    �7    �7    7    (7    P7    �7    �7    �7    �7    0     8     D6    t6    �7    �7    �7    �7    <7    \7    �7    �7    �7    �7    �7    �6    �7    �7    �7    �7    P7    p7    �7    �7    �7    �7     7     �6     �7     �7    !7    !7    !t7    !�7    !�7    " 7    "7    "7    "(7    "�6    #7    #7     c�h�w��4��]�S #$7    #47    #�7    #�7    #�7    $ 7    $(7    $87    $H7    $�6    % 7    %(7    %87    %H7    %�7    %�7    %�7    &47    &<7    &L7    &\7    &�6    '87    '@7    'P7    '`7    '�7    '�7    (7    (L7    (T7    (d7    (t7    (�     (�     (�6    ),6    )l7    )t7    )�7    )�7    )�7    *7    *<7    *�7    *�7    *�7    *�7    +86    +�7    +�7    +�7    +�7    ,7    ,(7    ,P7    ,�7    ,�7    ,�7    ,�7    -L6    -�7    -�7    -�7     d���]"��@� -�7    .7    .<7    .d7    .�7    .�7    .�7    .�7    /`6    /�7    /�7    /�7    /�7    0,7    0L7    0t7    0�7    0�7    0�7    0�7    1p6    1�7    1�7    1�7    1�7    2D7    2d7    2�7    2�7    2�7    2�7    2�7    4l6    4�     5x6    5�     5�     6 6    6�6    6�     76    7     7$     7@6    7L     7�     7�6    7�     7�     8(     8L6    8`     8h     8�7    8�7    8�7    8�7    9     9 6    9�6    9�     :7    :7    :7     e���e��	&��� :,7    :8     :@     :�7    :�7    :�7    ;(7    ;07    ;@7    ;P7    ;�6    <D7    <L7    <\7    <l7    <�7    <�7    =7    =X7    =`7    =p7    =�7    >6    >X7    >`7    >p7    >�7    >�7    ? 7    ?(7    ?l7    ?t7    ?�7    ?�7    @,6    @p7    @x7    @�7    @�7    @�7    A7    A@7    A�7    A�7    A�7    A�7    B      B(     B46    Bd6    B�7    B�7    B�7    B�7    C,7    CL7    Ct7    C�7    C�7    C�7    C�7    Dp6    D�7    D�7     f�}�S���}�SY D�7    D�7    E@7    E`7    E�7    E�7    E�7    E�7    E�7    F�6    F�7    F�7    F�7    F�7    GT7    Gt7    G�7    G�7    G�7    G�7    H7    H�6    H�7    H�7    I7    I7    I|7    I�7    I�7    J7    J7    J 7    J07    J�6    K7    K7    K 7    K07    K�7    K�7    K�7    L7    L$7    L47    LD7    L�6    M,7    M47    MD7    MT7    M�7    M�7    M�7    N@7    NH7    NX7    Nh7    N�6    O6    O$6         [�D ��       T   H  g�2�D�$���Š� �       '�    [�D3P                   (      �  ,(    �6     �6    �6    �6    t7    �7    �7    d     �6    �6    p6    x6    �6    L7    \7    �7    �7    7    L6    \7    l7    	     	<6    	P     	X     	�  	� 	�"    
@     
H          $     �6    �     D     H     X     p6    |     �     x     �     �     �     �     �                ,6    L     X6    �     �     �     �     �     �      h����J�ITQ�� �     �     �6         x     �6    �     �     �     �     \     l6    �6         T     x6    �     �     �7    �7    0     @6    �6    �     7    ,7    8     @     �7    �7    �7    ,6    <7    L7    �6    ,7    <7    �7    �7    �7    ,6    <7    L7    $6    ,6    �6    �6    �7    �7    �7    7    ,7    T7    �     46    �7    �7    �7    7    D7    �6    �7    �7    L6     i+QN��V#g� �7    �7     7     47     \7     �6     �7     �7    !D6    !�7    !�7    "7    ",7    "T7    "�6    "�7    "�7    #�7    #�7    #�7    %6    %6    &p6    &�6    &�6         [�D �`       T   H �       K�    [�D3�                   (     �  4     �      �      �      �      �      �          1               86    L     T     �     �     �     �     �1     �     �     �6    �#     6    �     �6    (6    �      j��_SQ%� �     �     �      6         06    <     �     �6    �     �          <6    P     X     �7    �7    �7    �7    �     6    �6    �     �7    �7    7    7    (     0     �7    �7    �7    7     7    07    @7    �6    	7    	 7    	07    	@7    	�7    	�7    	�7    
,7    
47    
D7    
T7    
�6    ,7    47    D7    T7    �7    �7    �7    @7    H7    X7    h7     6    H7    P7    `7     kROs<^oJ�Bp� p7    �7    �7    7    T7    \7    l7    |7    6    `7    h7    x7    �7    �7    7    07    l7    t7    �7    �7              0#     T6    �     �6    d6    �                46    <     H     d6    p     �6    �     �     6         $     t     �6    �     �     �7    �7    �7    7    T     l6    �6    $     P7    X7    h7    x7    �     �     �7    7    07    t7    |7     l�n�r�k3�=Do �7    �7    ,6    t7    |7    �7    �7    �7    7    D7    �7    �7    �7    �7    H6    �7    �7    �7    �7    7    47    \7    �7    �7    �7    �7    d     l     t     |     �     �1     �     �     �6    �#     �6    �     �6    6    �     �     �     �     �6    �     6         h     �6    �     �     �      6     0      8      d7     l7     |7     �7     �      �6    !h6    !�      m.7á���=4$ !�7    !�7    !�7    !�7    "     "     "l7    "�7    "�7    "�7    # 7    #7    # 7    #�6    #�7    $ 7    $7    $ 7    $�7    $�7    $�7    %7    %7    %$7    %47    %�     %�6    &�     &�6    '6    '�     '�     '�     '�6    '�     '�     (6    (     (46    (@     (�     (�6    (�     (�     )     )@6    )T     )\     )�7    )�7    )�7    )�7    )�     *6    *�6    *�     *�7    + 7    +7    + 7    +,     +4     +�7    +�7     ni�-V�F��{� +�7    ,7    ,$7    ,47    ,D7    ,�6    -7    -$7    -47    -D7    -�7    -�7    -�7    .07    .87    .H7    .X7    .�6    /47    /<7    /L7    /\7    /�7    /�7    07    0H7    0P7    0`7    0p7    0�     0�     16    1\7    1d7    1t7    1�7    1�7    27    2,7    2p7    2x7    2�7    2�7    3#     3<6    3�     3�6    4L6    4�     4�     4�     56    5     5(     5D6    5P     5t6    5�     5�     5�6    6     6     6\     6�6     oN(~0���c��ߩ 6�     6�     6�7    6�7    6�7    6�7    7<     7T6    7�6    8     887    8@7    8P7    8`7    8l     8t     8�7    8�7    97    9\7    9d7    9t7    9�7    :#     :(6    :�     :�6    ;86    ;�     ;�     ;�     < 6    <     <     <06    <<     <\     <�6    =,     =H6    =�6    >@     >T     >X     >p6    >|     >�     >�6    >�     >�6    >�     ?,     ?P6    ?d     ?l     ?�     ?�6    ?�     ?�     @(7    @07    @@7    @P7    @�      p$Q7�Pl�fCw� @�6    A,6    Al     A�7    A�7    A�7    A�7    A�     A�     B07    BP7    Bx7    B�7    B�7    B�7    B�7    Cd#     C�6    D     D06    D�6    E      E4     E8     EP     Ep6    E|     E�6    E�     E�     F6    F0     F8     F�     F�6    F�     F�     F�7    F�7    G7    G7    Gh     G�6    G�6    H8     Hd7    Hl7    H|7    H�7    H�     H�     H�7    I7    ID7    I�7    I�7    I�7    I�7    J0     J�6    J�6    K6         [�D�  q,P�E-s��       T   H �        h    [�D4p                   (      �  4     �6     7    7    7    (7    �7    �7    �7    7    7    ,7    <7    �     �     �6    ,7    47    D7    T7    �7    �7    �7    @7    H7    X7    h7     6    D7    L7    \7    l7    �7    �7    7    P7    X7    h7    x7    �     �     0     8     @     H     T     X1     `     l     �6    �#     �6    P     l6    �6     rH"-��� ����- 	\     	p     	t     	�     	�6    	�     	�6    	�     
4     
X6    
l     
t     
�     
�6    
�          07    87    H7    X7    �     �6    46    t     �7    �7    �7    �7    �     �     87    X7    �7    �7    �7    �7    �7    x     �6    H     d6    �6    \     p     t     �     �6    �          (6    <     D     �     �6    �     �      7    7    7    (7    t     �6    6    D      s�0Ek���%���� p7    x7    �7    �7    �     �     7    (7    P7    �7    �7    �7    �7    T6    �7    �7    �7    �7     7    @7    h7    �7    �7    �7    �7    `6    x6    �6         [�D+        T   H �        +�    [�D5                    (      �  4     �      �      �6     �6     7    (7    87    H7    �7    �7    �7    47    <7    L7    \7    �6    47    <7    L7    \7    �7    �7    7    H7     t�Wj�A�n� P7    `7    p7    6    T7    \7    l7    |7    �7    �7    $7    h7    p7    �7    �7    #     46    �     �6    D6    �     �     �     	6    	$     	0     	L6    	X     	�     	�6    	�     	�     
4     
X6    
l     
t     
�7    
�7    
�7    
�7         ,6    �6    �     7    7    (7    87    D     L     �7    �7    �7    47    <7    L7    \7    �#      6    �     �6    6    �     �      u��(���>l.D �     �6               (6    4     X#     x6    �     6    �6                    86    D     P     l6    x     �6    �     �     6    $     ,     |     �6    �     �     �7    �7     7    7    \     t6    �6    ,     X7    `7    p7    �7    �     �     �7    7    87    |7    �7    �7    �7    <6    �7    �7    �7    �7    7    (7    P7    �7    �7    �7    �7    |  x �"     vz�+�`nAU�8B (     0     �6    �7    �7    7    7    |7    �7    �7    7    7     7    07    �     �     �     �1     �          $6    8#     \6    �     6    l6    �               46    <     H     d6    p     �     �6    �     �      L      p6     �      �      �7     �7     �7     �7    !,     !D6    !�6    !�     "(7    "07    "@7    "P7    "\     "d     "�7    "�7    #7    #L7    #T7    #d7    #t7    $6     w"��9M��<x�> $T7    $\7    $l7    $|7    $�7    $�7    %$7    %h7    %p7    %�7    %�7    & 6    &h7    &p7    &�7    &�7    &�7    '7    '87    '|7    '�7    '�7    '�7    (<6    (�7    (�7    (�7    (�7    )7    )(7    )P7    )�7    )�7    )�7    )�7    *H6    *`6    *x6         [�DV�       T   H �        �    [�D5�                   (      �  4     �      �      �6    7    7    ,7    <7    �7    �7    �7    (7    07    @7    P7     x�?1���aA# �     6    �     �6    6    �     �     �     �6    �     �     6          l     �6    �     �     �      6    4     <     h7    p7    �7    �7    �     �6    l6    �     �7    �7    �7     7              p7    �7    �7    �7    	7    	7    	$7    	�6    
$     
H6    
\     
d     
�7    
�7    
�7    
�7         6    �6    �      7    7    7    (7    4     <     �7    �7    �7     y����R���� $7    ,7    <7    L7       ("    �     �                     $1     ,     8     T6    t#     x#     h6    �     �     �6    X6    �     �     �6    �     6    $     p     �6    �     �           $6    8     @     l7    t7    �7    �7    �     �6    p6    �     �7    �7    �7    7              t7    �7    �7     7    7    7    (7    �6    �6    �6         [�Dn�       T   H  z��+/V/�&���` �           [�D6                    (      �  4     �6     7    7    7    (7    �7    �7    �7    7    7    ,7    <7    �6    7    7    ,7    <7    �7    �7    �7    (7    07    @7    P7    �     6    �     �6    $6    �     �     �     �6    �          $6    0     |     �6    �     �          06    D     L     x7    �7    �7    �7    �     	6    	|6    	�     	�7    	�7    
 7     {݅+/\N"(�j 
7    
     
$     
�7    
�7    
�7    7    7    $7    47    �6    7    7    $7    47    �7    �7    �7     7    (7    87    H7    �6     7    (7    87    H7    �7    �7    �7    47    <7    L7    \7    �6    47    <7    L7    \7    �7    �7    7    H7    P7    `7    p7     6    L7    T7    d7    t7    �7    �7    7    `7    h7    x7    �7    46    �     �6    H6    �     �      |�p�o�Ӈ�D�� �            6    ,     x     �6    �     �          ,6    @     H     t7    |7    �7    �7    �      6    x6    �     �7    �7    �7    7               |7    �7    �7    7    7     7    07    �6    7    7    7    ,7    �7    �7    �7    7     7    07    @7    �6    �6    �6         [�D��       T   H �        �    [�D6�                   (        4     �     7    $7    L7     }�p��řZ<��� x7    �7    �7    <7    L7    \7    �6    $6    X6    �6    �6    $7    D7    l7    �6    �6    �6         [�D��       T   H �       �    [�D7@                   (        ,�   �6     �6    6    �6    �6    �7    �  � �"    \     d     |     �               �6         <6    P     X     �#     �     L6    T6    	|7    
X7     6    6    06         [�D��       T   H �        	�    [�D7�  ~x?���9�6�                   (      $  4     �7    7    T7    \7    �6    �           6    �6    �          (6    4     `     �7    �7    7    T7    $6    <     `6    �     �     �     \     �6    �     �     �7    �7    �7     7    �6    �6    �6         [�D�0       T   H �       8    [�D8`                   (        4    �     �     $     <6    �6    �     <6    D     P     l6    x     �6     ���aѕ�_�ua/ �     <     h6    |     �     �     <6    �6    �6    d6    l6    	87    
6    
,6    
D6         [�D��       T   H �       #0    [�D8�                   (      Z  ,      "    #     p#     |6    �6    �6    T7    x7    <  8 P"    d  ` x"    �  � "    h6    �  � �"    	6    	 6    	�  	� 	�"    
7    
87    
`7    x7    �7    �7    �6    �7    �7     7    �7    �7    T     �6    t7     �ǀ�.^'S��"�� �7    �7    7    $7    L7    47    T7    |7    d7    �7    �7    �7    �7    �7    �7    �7    7    06    86    �6    <     D     �  � �"       � "    x     �  � �"    �6    �6    @6    H6    h6    �6    �6    �6    �6    T7    �7    �  � �"    �  � �"     6     6    !P  !L !d"    !|6    !�6    "�  "� "�"         [�D��       T   H �        �    [�D:                   (        , @   ��"�p��4�Q<�      [�D         T   H �       �    [�D:�                   ,        0@  7    T7    87         [�D-�       T   H �         �    [�D9�                   0        4             �                   �        "      "�  
        �x     -   �        ۸     F�  8        ވ     N   P`        ߸     ��  '�        ��     �`  L         ��    �  x        �    +   +�        �    V�  �        0    n�           �    ��  ��b�7�Z	�          �    ��  �        �    ��  	�        �    �0  H        @    ��  #@        x    ��   �        !�    -�   �        "x          D 	�               L �               P $               L PP        ,       D T � 	� 	� 
%X %� '�               L K�               L h               L � � 
+�               L ( , 
�               L                L �               D � � 
�               L   �=��-��yZqzF	�               L 4          B    D    � @ � P "T #x "| #� "� + " #� "� #	d "	� +	� "	� #
T "
� 5� "( 5 "� 5� "T 5@ "� 5p "� 5� "� 5� " 5  "D 5\ "� =� "� # " #  "� E� F� E� N� O� N� O� N | E � X!, E!H a!d E!h F!p E!� f"D g"� f"� m# f#,               @  �               L � r      �      s                                                                                                                 �O���������                                                  	   
                                                                                                                                                                                                        0                         �    � @               E     �  �    � @               C     �  �    � @               A     �  �                        @     �    ��9�IW���=U    � @                       U    � @               ?        �    � @               =       �    � @               ;     �  �    � @               9       U    � @               7 f      �    0 �               5       �    � @               3     �  �    � @               1     �  �    � @               /     �  �    �                       �                                      �                                  ����&}s_�o��                                                }                      ����                                        � �                         -     �                                   @ �� �                       -     �                                   @ �� K                       +                                 ��������                �a�8���@���H���P���X|�� (�!��`\  �A  < D� 3�  | �A݀`}  �|  c~  �~�- @� ;`  �~�H  $;��cc  c�  K���;`  �~;` �~  �?�'��"���A݁�8!@� (|��a�;N� !    ����[�D"x          H  �        @           [�D/    ��                                         w��� (w��� *w��� �0w��� �w��� ��w����w�����w����`w��� �                        �  ��                         [�D  [�D �        [�DC�4�� 54�� 7�        [�D.�4�� 1`[�DD@[�DE�        [�D1 4��  [�D)@[�D'h                                �       =      �   F �    [�D0         ��,+����                        u�N��  �4 9�_�3١        [�DGP[�D;0                                                                                                                                                                                                                                          
0                  
    [�D "�[�D/ [�D "�[�D$�4��   4�� .Pw���                                     �   �  v                      .�;       �    [�D - [�D/ [�D - [�D$�4��  `4�� .�w���  �                          ��о�kD�j�/�          `   ;  -                      �K�       8    [�D F�[�D/ [�D F�[�D$�4�� !84�� .�w���  �                                  �   �  �                      �th�       P`    [�D N [�D/ [�D N [�D$�4�� !x4�� / w���  �                                  �   �  �                      �ս@       '�    [�D ��[�D/ [�D ��[�D% 4�� $4�� /Hw��� 8                                  �    �                      ���       L     [�D �`[�D/   �!������y��[�D �`[�D%04�� %P4�� /�w��� �                                  �   �  x                      �       x    [�D�[�D/ [�D�[�D%H4�� '�4�� /�w��� �                                  @   I  5                      �w��       +�    [�D+ [�D/ [�D+ [�D%`4�� (�4�� /�w���                                   �    �                      ���       �    [�DV�[�D/ [�DV�[�D%�4�� )�4�� 0(w��� X                                     <  ��S�M�V�sy3W  �      	                l8            [�Dn�[�D/ [�Dn�[�D%�4�� *�4�� 0Pw��� �                                  `  ,  �      
                ���           [�D��[�D/ [�D��[�D%�4�� +�4�� 0xw��� �                                  �   +  *                      �V�� @     �    [�D��[�D/ [�D��[�D%�4�� , 4�� 0�w��� �                                  `   m  H                      ��0 @     	�    [�D��[�D/ [�D��[�D%�  ����H�w�� �4�� ,h4�� 0�w���                                   �   T  C                      ��L�       H    [�D�0[�D/ [�D�0[�D&4�� ,�4�� 0�w��� @                                      �  w                      |�e�       #@    [�D��[�D/ [�D��[�D& 4�� - 4�� 1 w��� p                                  @                           �: �      �    [�D-�[�D/ [�D-�[�D.(                                                          @  O  �            �Pԩ�N���j�            ��A        �    [�D��[�D/ [�D��[�D'8                                                          `  +                         oPg�       �    [�D  [�D/ [�D  [�D'P                                                             =                         ޻��  �                         @[�D�x                                                                   �                 �[�D۸                                                                 �     �'��/2�O�=!              0[�Dވ                                                                 �                 ([�D߸                                                                 �                  �[�D��                                                                  (                  ([�D��                                                                 j�                 �[�D�                                                                 *@                 P[�D�          ��{,
B���=>                                                         B@                 �[�D0                                                                 &@                 �[�D�                                                                 6@                 [�D�                                                                 �                 @[�D�                                                                  �                 x[�D�                                          ���^���⛷d`                                           8[�D@                                                                 @                 ([�Dx                                                                      
               `[�D"x                                                                                      `[�D!�                                                                   @                   x[�D"                                                                   @     �)��9�k�qT��   	                          "   &      3                  [�D �                [�D p                        [�D �[�D �[�D  [�D �                                        [�D`��HY3m�    C                                                                                                                                                               �   �   w���Ր        w���א        w����P                         000`p00 
 %��������@@@@@@@@@@@@@@@@@@@@@@�����@@@@@@@@@  ��T�C0�����?K@@@@@@@@@@@@@@@@                  0                            `                 �     	�      �     
$      �     �                 `   	  4      �   	  �      H     �      h     D      �     \           �      0     �      H     �      `     \      x           �     8      �     `      �     |      
           
0     "�      
H     #      
�     "�  �                 �             �             �                                    ���e�Ǐ1(�
                    h   	          x   	          �   	          P             `             p                                                      8             P             h             �             �             �             �             
              
8             
P             
�         0   �              d             p            �            �                        �            �             t            �             p         ���UOL}1I�i%j     X            h            �            �            \            �            �            �            �                                     "<            $\            &p            (�            *�            ,�            .�            0�            3            ;d            =�            ?�            A�            C�            F            H            JD            LX            N|             d            �         ��=}8=��C�)Kh     �            �            �            �            `            `            ,            �                        T            �            �             �            "�            $H             p            T            
h            |            �            �            �            �            �            #4            %H            ,X            .l            0�            2�            9�            B�         ��"zx�+_��A     I�             p            P            |            �                         �            �             p            p            �            �            p            �            �            D            #�            %�            '�            )�          	   p          	  d          	  	8          	  `          	  <          
   p          
  P          
  d          
  H          
  \          
  p          
  �         ��d��ASN>��^    
  �          
  D          
  T             p            $            8             d             p             p            �            	|            
�            $            �            P            �            �            �   	            
         @            �            !D             l            `                                                                                                                                         ��s"r@���Րբ "  �  [�D        4��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ��rO�G�)s �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��s�Xo   s@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   s`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   s�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   s�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   s�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   s�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   t                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ��s�Xo   t                \���� @]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@%\�����������LL% \������������ @�\������������ �@\�����������nn% \������ ���������@  \��������   �����   �����M]@������K@������M]@������K@   �M] \������ Ù���Ƣ���  ]}% ����M]@������K@ Ù���Ƣ���  @�@�����������  ��% �����M]@������K@���������@  a��@l���`�K�%   @� lBFw�%     
�        
`            �          �   a㉣��@M     K            �         �����s��X�V�aÙ������ā��@M�z   @� aי������@M�������@��K�@M����@���Ö���k@����]]%   @�� ������% a㨗�@aÁ�����% aׁ���@�@�@�%   a㨗�@aƖ��%��% Ö����� a⤂����@a㨗��%aՁ��@a��%  @�% a��Ɩ��@a @z@ aŕ������@a払����ŕ������% ��� @@aƖ��@LL@a��@�@�@�@nn%@@aי��Ⅳ@�@a���@aㅧ�@�%      ����������      �����������     ���������@�����������������@@@@@@@@     �����   ���������@�����������������@@@@@@@@     �����   [�D �X[�D ��  �    [�D ��[�D ��[�D ��  �    ���������@�����������������@@@@@@@@     ��������  ��0~���`���������������������@@@@@@@@     ����������      @�@���  a㨗�@aׁ��%    aׁ����@�@�@�%  aم�������@�@�@�%       aÖ������@      aӅ����@������% �@�@�@�@���������@      ���������%      �������@@@      a㨗�@aׁ���%   aÖ���@ aԅ����@�@�@�@a҉��@� [�DD�[�D+   e    [�D+ [�DE[�D+   e    ��������������  ����%   ����������@�����@�@%    [�Dd�[�DV�  �    [�DV�[�DeL[�DV�  �    @�����@�@       ���������@      a≩�@  aٖ��@�@�@�%    aɕ��@�@�@�%    ���������%      ll���%  ��������  ���dza;��Y�<��      ������������    Ó���Ƣ���      ����������      ������������    [�D��[�D��  �    [�D��[�D�[�D��  �    ����������      �����������     �@���������� ����������      ������� ř���@  �������@@@����  \������ ���������@      [�D��[�D��        [�D��[�D�|[�D��        [�D�$[�D��        [�D�4[�D��   �    [�D��[�D�� BA    [�D��[�D�� BA    ���������@      [�D��[�D��   �    �����   �����   [�D��[�D��   �    [�D��[�D��   �    @@@@@@@@  �|mMp�&���@@@@@@@@@@@@@@@@@@@@@@@@��������@@@@@@@@@@@@@@@@@@@@@@          P      @@       �        �����  ������������    �@@@@@@@@@@@@@�@@@@��������@@����������\����@@@\����@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�����������������������������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����������������������@@@@�������@@@��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �`v�<�zx���w@@@@@@@@@@@@@@@@@@@@@@@@[�D��[�D�� BA    [�D�8[�D��   �    [�Dٔ[�D�� BB    ���������������@@@@@@@@@@@@@@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����������@@@@�����������\����@@@\����@@@@@@@@@@@     [�D�X[�D��   �                                                                                                                                                                                                                                                                                     �w��8��L~*                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��s�Xo   u     \         K    P     �   @U     
��    
�� UX ��           �� (   � � � �         �             
                                   �                            (             @               P         �                  P                              �                          �        @                                    @@                P  �     �  �    
                                A                                @                                               ���iK7��T&�                                                                       �                                               �                                                                               @@                                               �                                                                                              �                                @                                               @                                �                                  �����8-2�
�       $  D         	�    P                   �                            @�                        �                       �                        T                                                                     
                    ��                                            *�          T                   l     d  �    
    �    @                       �                                             @                                               @�                        �#�s�t���                                               �                   @                       �                                             @                         @                                                              �                                         @                                                                         @                                                                                  �               �         �    
                                           ��3��X���=�        @                                                                                                                            @       d         
�    
                                �                �                                                                                               @                                                     �                 �                                                        P                �                                        �     �	{�:��� j�'�      �    
                �                       @                                                                                                                                 �     �         -    
                                �                                                     @                                               �                                                                   �                    H         �    
                                                  ��w�EЃ ��`   h         �    P                                            
                                     T             
           �                                                         `             
         �                         �  T                                ,         �                                                                !           �                    �                                                                         @                            ��r��0�V`�                                                                                  ]          E   �   		
 !!"#$%&'())*+,-./011234567889:;<=?@ABE      .               
"#$'()-                  D      E          -  g    !$%&'()*+,,-./01236789:;<?      F          .  �    !"#$%%&()+,./0122344567899;<<>A     :          "  �   
 "#$'*+.03469         %            ,   
      -     �J�/���n�p�m         K   
 "#$'      %            v         %            �   	                  �   	                  �   *,-.025                   	       (                !"$(   X             �    A�                  
                         A�          �               \�����m�������   �����   ������������   
����������   �������   
����������   mm�����   �����������   ����   \�����m��������   \����  �5��|د����S�m��������   	���������   	���������   	���������   ��������   ������   �����   	���������   �����������   
����������   ��������������   ������������   	���������   	\����m���   \�����m�������   m����m����m���   m����m��m���   m����m���m�����m���   m����m����m��   
m����m����   m����m����m����   
m����m����   m����m�����m��   m����m�����   
m����m��m�   ��������   m����m����m�   m����m������m����   
m����m����   m����m������   m����m�m������m�   m����m�m��m�   m����m�m�����m�   m����m  �=�"\P?�R��>����m�����   m����m����m��m�   m����m����m��m�   m����m����m����m�   m����m��m���m��   m����m��m����   m����m����m�   m����m���m���m�   m����m����m���   m����m���m��������   �@��@��ą�����ň   �@��@���È   �@��@������������ɕ��   �@��@���ŗ����            4�� 5x4�� 7�                                                4�� 7�                                0   "          )   "   �     D   b   �     W   |   �     {   �   �     �   �   �     �   �   	�     �  h   �     �  z  ��u!�u���b�E   �       �   �       �   E        �   �       �   �       �   �       �   C        �   �     l     �     �     A      �  ,   �     �  A   !�     �  _   ?      �  s   =      �  �   ;      �  �   #�     �  �   9      �  �   7      �  �   5      �  �   3      �  �   %�     �     1      �     /      �  S   -      @  g   +      D  w   '�     G  �   )�                                                          4�� 8h4�� 8�          �!�����0��4�� 9�                        4�� 8�                        ����$�t  +�                             h             +�      	                                                                                                         �   	             X      �             `  h  @             	�    �             
�   �  �             �     P                �  �                  �                 0  *�             R     +r           �                �  �         p  ���V�.I��v�$  p         �  �         �  �         �  �         �  �         �           �  @         �            �   �         �  )`                                                                                                                                                                                                                                                                                                                                                                              �i�A���4 t֋                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��s�Xo   v�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   w   ��  [�D                   e                  E   �   		
 !!"#$%&'())*+,-./011234567889:;<=?@ABE      6                       
"#$'()-     (                    D      M                  -  g    !$%&'()*+,,-./01236789:;<?      \      P           /  �    !"#$%%&&()+,./0122344567899;<<>A                 B                  "  �   
 "#$'*+.03469         -                    ,     ���ZrI���ř��
      D      8             K   
  "#$'                  -                    v         -                    �   	      &                    �   	     8      ,           	  �   *,-..025               $                        	       0                        !"$(   `                     �    A�                  
                         A�  $8     �     �                d        ��f!��u8�^!�          e                f                g                h                i                o               �                 p             !   q             "   r             #   t             $  �             %   x             &   |             '   �             (   �             *  �             +  p             ,  �             -  �             .  �             /  @             0               1               2  �             3  �  ���I}$x|�d�             4                5               6   �             7   �             8   �             9   �             :   �             ;   �             <                =  0             >  @             ?  P             @  p             A  �             B   �             C   �             D   �             E   �             F   �             G  �             H  P             I  `             J  p             K  �             L  �            ��'t�<v�M[   M  �             N  �             O  �             P   �             Q   �             R   �             S   �             T   �             U   �             V   �             W                �  �             �  !             �                 �  �             �                �   P       w   �   @       w      0       w             w             5                 �               �            �               �    ���P�o���Ɵ/          �            	   �          
                  �                           �                            �            0               �            @               �            P               p            `               `            p               P            �               @            �               0            �                             �            #  �5��lt�����&               $  �       �  %           �  &  �       �  '  �       �  +   �            , �       �  . �     �  �  /  �     �  �  0 @     �  x  1 �     �  5  2 �     �  �  3 �     �  �  4 �     �  �  6  �          7 0     �  -  8  �     �  �  9  �     �  *  : �     �  w  <        C  =         H  >   �            ?   �            @ �     e  -  A  �            E �       � !6c��c�f(�  �  F �       �  G @       w  I  �    x  H  J               K          �  L  	             M  �            N         H  O          H  S              T              U              V              X              Y              Z  %p            [              ^          �  b              k         d  -  o  	�            p  �            r  �       �  s  �       �  t              u     ���$u{*9�JP�x            y �       5  | 0       x  }  
0            ~          H            H  �         d  �  �  $            �  &            �  (            �  ,            �  0            �  $       H  �  �            �  �            �  )`            �  0            �  �            �  �            �  �            �               �  P            �  p            �              �  �            �  �            �M�l���1oդ  �               �  �            �  �            �  0            �              �  0            �  @            �  P            �  `            �  p            �  �            �  �            �  �            �  �            �  �            �  �            �  �            �  �            �               �              �               �  0            �  @            �  P            �  `            �  p     �k��i�+'o'         �  �            �  �            �  �            �  P            �  �            �  @            �  P            �  �            �               �  �            �               �   0     �  v  �           v  �           v  �          v  �  �            �       �  -  �  p       -  �           -  �  �       -  �       ��  -  �         -  �          -  � �     0  -  �  �     �  -  �  ��>�fEX�vK  0       -  �  @       -  �  P     
  -  �        -  �  `       -  �  �            �      �  �  � �     0  �  �        �  �  �        ��  �  �  �            � @     �  �  � �       �  �  �       �  � �     0  �  �         
  �  �          �  �           �  �   0       �      @    ��  �   �       �    @       �   �       �    P       �    `       �    p       �W��@���Xxޮ  �    �            	        �  �  
  p              �     0  �    `       �    `       �             �    p       �            �             �     0      �    �       �    @       �    P       �     �            ! 4       x  " �     �  x  #                $           x  %          x  &           x  '  �       x  (   0       x  )   @    ��  x  *  @       x  +  �  �u3M�~�x�9cK       x  ,  �       x  - �       x  . @     0  x  / �       x  0 �       x  1  P       x  2  p       x  3 �       x  4 �       x  5         x  6        x  7         x  9  �            : `     �  5  ;  �       5  < �     0  5  =           5  >          5  ?           5  @ �       5  A   0       5  B   @    ��  5  C  @       5  D �       5  E �       5  Ƽ�����_`�  F  P       5  G  p       5  H �       5  J  �            K `     �  �  L �       �  M  P       �  N �     0  �  O           �  P          �  Q           �  R P       �  S   0       �  T   @    ��  �  U  @       �  V `       �  W p       �  X �       �  Y �       �  Z �       �  [ �       �  ]  �            ^ P     �  �  _  �       �  ` �     0  �  a        ǧ=���LEՄ�(�     �  b           �  c   0       �  d �       �  e   P       �  f   `    ��  �  g  `       �  h �       �  i �       �  j �       �  k  p     
  �  n  �            o `     �  �  p �       �  q  �       �  r �     0  �  s           �  t           �  u   0       �  v �       �  w   P       �  x   `    ��  �  y  `       �  z �       �  { �       �  |  p     
  �  }  ���ҧ.+|0|�  �       �  ~ �       �  �  �            � P     �  *  �  �       *  � �     0  *  �        �  *  �        ��  *  �        
  *  �  �       *  �         *  �  �            �  %       H  �        �  H  �  0       H  �           H  �        
  H  �   �       H  �   �       H  �  �     0  H  �   �       H  �          H  �           H  �   0       H  �   @       H  �   P       �R=��Po�r��  H  �   `       H  �   p       H  �   �       H  �   �       H  �   �       H  �   �       H  �  �            �         C  �       �  C  � �     0  C  �         
  C  �          C  �  `       C  �           C  �  p       C  �   0    ��  C  �  0       C  �  @       C  �  P       C  �  �     �  C  �  �            � `     �  w  �           w  �  �       w  �          w  �      �l�1zs���n�       w  �  �       w  �   0    ��  w  �  0       w  �  @       w  �  �       w  �  P       w  �  �     �  w  �  `       w  �  p       w  � �     0  w  �   (            �  P            �  `            �  p            �  �            �              �             �             �  0     d     �  �            �  �            �  �            �   0            �   @            �           �  ��S��nbx[�I�  �   P            �  �            �   `            �  �              @       H    P       H    `       H    p       H    �       H    �       H    �       H    �       H    �       H    �       H    �       H    �       H   P       w   `       w   p       w   �       w    �       w  ! �       w  " �       w  # �       w  $ �       w  ?        ���Ã���V�Q                      ��������@@@@@@@@@@@@@@@@@@@@@@�        �                                                               �                                                   I ��                           %00         
                                                                                                                                                                                                                                                                                       ͩ�\]���                  �     H����                                           u  Y            0           T                                                                                                                                                                                                                                                                                                                                                                                                   ����R����p                            	 H                        	 H                         H                                                                                                	                   p � �                                                                                     p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p �   ��<�*T5�m��<�  	                   p � �                     p � �                     p � �                     p � �                     p � �  	                   p � �                     p � �                     p � �                     p � �                     p � �                                             �   =    x � �                     � � �                      � � �              �        � � �             0        � �   Б����!iP��<�              �        � � �              @        � � �                    p �                        � �                      � �  	                   p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p � �  	                   p � �  	                   p � �  	                   p �   ѕZsr��drbX%��                      p � �                      p � �                      p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p �   ҕ|���8�8Q܀              H       p � �                     p � �                     p � �              
       p � �                     p � �                     p � �              
       p � �                     p � �              �   P    x � �                                                                                                                                                                                                                                Ӑy��	�i�6�0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ԉs�Xo   z�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   Չs�Xo   z�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ։s�Xo   z�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ׉s�Xo   z�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ؉s�Xo   {                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ىs�Xo   {                                                                                                                                                                           W   m      P    x @ �                                                                                                                                                                                                                                                                                                                                 ڈ��Do  �"�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ۉs�Xo   {`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ܉s�Xo   {�                                                                                                                                                                                                                                                                                                                                          W      c   P    x @ �                                                       ` � �                      ` � �                      � �  	   w              � �   ݉vR�����̀  	   w              � � �  	   w              � � �  	   w              � � �  	   5              � � �  	                  � � �  	                   � � �  	                  � � �  	                   � � �  	                  � � �  	                   � � �  	                  � � �  	               	    � � �  	                  � � �  	               
    � � �  	                  � � �  	                   � �   ޕ�ҵ:�D� C܀  	                  � � �  	                   � � �  	                  � � �  	                   � � �  	                  � � �  	                   � � �  	                  � � �  	                   � � �  	                  � � �  	                   � � �  	                  � � �  	                   � � �  	                  � � �  	                   � � �  	                  � � �  	                   � �   ߕ���:� ���{��  	                  � � �  	                   � � �                                                                                 f    p � �      �              p � �     �              p � �     �              ` � �     �              p � �                                                             `                               ` � �     �              p � �          /  O               �       �       p �   ��荶h4X���+��     �       �       p � �     x       �       p � �     5       �       p � �     �       �       p � �     �       �       p � �     �       �        p � �          "  �                          ]    ` � �     -       �   !    p � �     �       �   "    p � �     *       �   #    p � �     w       �   $    p � �                      `   �  	   C          %    � � �     H          &    p � �                 '    p �   �̄df�r���)�                 (    ` � �     -       e   )    p � �                 *    p � �                      `   �            �      �                            	 H   �          +    p � �     �          ,    p � �     w          -    p � �            b              H      x   .    p � �                 /    ` � �     �              ` � �              �   0    p � �             �   1    p � �     H          2    p �   �����׆fm��     H          3    p � �               �       `   �                      `   �               
       `   �                 4    ` � �                 5    ` � �                 6    ` � �                 7    ` � �                          8               8    ` � �                 9    ` � �             �   :    p � �                 ;    ` � �                      `   �                      `   �     �          <    p �   �!>�U��hG���               
       `   �                      `   �               
       `   �                 >    ` � �               
       `   �                      `   �                      `   �                      `   �                      `   �                      `   �                      `   �               d       `   �     -       d       p � �                      `   �                      `   �                            �><��'����)P             \   ?    p � �                 @    p � �                              �          A    ` � �     �          B    ` � �                 C    ` � �                 D    ` � �          %  y                      E                    ^  �              5          E    ` � �                      `   �                         	    x          F    ` � �                 G    p � �     H          H    p �   �i㶢�/{IC/@�     H          I    p � �     �       d       p � �                 J    ` � �                                         K    ` � �                                    \                    Z  �                    \  �                    =  �                    &  j                    *  �                                     H               L    ` � �                 M    ` � �                 N    ` �   ��˵.~A�@�<�     H          O    p � �  	                    x � �                      x � �             �       � � �              P        x � �              �        � � �  	               �    p � �              �   �    p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p � �                     p �   ��Se{w���D��                     p � �                     ` � �                     ` � �                     ` � �                                              
       ` � �                                              
       ` � �                                              
       ` � �                                              
       ` � �                                              
       ` � �                                              
       ` �   �5&���|*��                                              
       ` � �                                              
       ` � �                                              
       ` � �                                              
       ` � �                                              
       ` � �                                              
       ` � �                                              
       ` � �                                              
       ` �   �v���nD:�L�                                              
       ` � �                                              
       ` � �                                              
       ` � �                                              
       ` � �                                              
       ` � �                                              
       ` � �                                              
       ` � �                 g    h � �                 h    h �   �v�(�m�k�QL�              �       p � �              �       ` � �                     ` � �                           0                         0                    � � �              
       ` � �                      ` � �                                                       ` � �                 Q    p � �     v       �        � � �     v          ^    p �    	   v          �    p �       v          R    p �                                  �T��}1��R|VP                        ` � �     -       �        � � �  	   -          �    p �       -          k    p �    	   -          �    p �       -      ��   �    p �       -          l    p �       -          m    p �       -       0        � � �     -       �   �    � �       -          _    p �       -          S    p �       -       
   �    p �       -          �    � �       -          �    p �                                  �]�hA��zt@                        ` � �     �       �        � � �     �       0        � � �     �       �   �    � �       �      ��   �    p �                                                        ` � �     �       �        � � �     �               � � �     �          �    � �       �       0        � � �     �       
   �    p �                                �          �    p �                                �          �    p �   �9�b5���b`�      �          �    p �       �      ��   �    p �    	   �          �    p �       �          n    p �    	   �          �    p �       �          o    p �       �          `    p �       �          T    p �                                                        ` � �     �       �        � � �              0   �    p � �                            �         /     �                                                              �+�?n0f�                              �       0        � � �     �          �    � �    	   �          �    p �       �          p    p �       �          �    p �       �          a    p �       �          q    p �                               �         �    p �    	   �          �    p �       �          b    p �       �          r    p �     �         /     �                                                              �Nz;��MQ�lee                                                     ` � �     x               ` � �     x       �        � � �                 c    p � �     x          �    p �       x          s    p �       x          �    p �    	   x          �    p �       x          U    p �       x      ��   �    p �       x          t    p �    	   x          �    p �       x          �    � �    	   x          �    p �       x       0        � �   �I���؜��  	   x          �    p �    	   x          �    p �       x          �    p �       x          �    p �    	   x          �    p �    	   x          �    p �    	   x          �    p �    	   x          �    p �    	   x          �    p �                                                        ` � �     5       �        � � �     5          �    � �       5       0        � � �     5          �    p �       5          u    p �   ��o��J��!�      5          �    p �    	   5          �    p �       5          V    p �       5      ��   �    p �       5          v    p �    	   5          �    p �    	   5          �    p �       5          �    p �       5          �    p �    	   5          �    p �                                                        ` � �     �       �        � � �     �               � � �     �          �    � �       �       0        � �   �����p8�ˉ�     �          �    p �       �          w    p �       �          �    p �    	   �          �    p �       �          W    p �       �      ��   �    p �       �          x    p �    	   �          �    p �    	   �          �    p �    	   �          �    p �    	   �          �    p �       �          �    p �    	   �          �    p �                                                        ` � �     �       �        � �   ��Ym�p�U1I�     �          �    � �       �       0        � � �     �          �    p �       �          y    p �       �          �    p �    	   �          �    p �       �          X    p �       �      ��   �    p �       �          z    p �    	   �          �    p �    	   �          �    p �       �          �    p �       �       
   �    p �                                                                                  ` �   �9-	֒� �3���     �       �        � � �     �               � � �     �          �    � �       �       0        � � �     �          �    p �       �          {    p �       �          �    p �    	   �          �    p �       �          Y    p �       �      ��   �    p �       �          |    p �    	   �          �    p �    	   �          �    p �       �       
   �    p �       �          �    p �    	   �          �    p �   ���}�Ұ8���                                                       ` � �     *       �        � � �     *               � � �     *       0        � � �     *       �   �    � �       *      ��   �    p �       *       
   �    p �       *          �    � �       *          �    p �                                                        ` � �     H               ` � �     H       �        � � �     H               � � �     H          �    p �   ��9���W�Wi���      H       
   �    p �       H          �    � �       H          �    � �       H       0        � � �                            H   H          �    p �    	   H          �    p �       H          d    p �       H          }    p �       H          ~    p �       H              p �       H          �    p �       H          �    p �       H          �    p �       H          �    p �       H          �    p �   ����}�_8��B�      H          �    p �                                                        ` � �     C               ` � �     C       �        � � �     C       0        � � �     C       
   �    p �       C       
   �    p �                              H	   C          �    p �       C          �    p �    	   C          �    p �       C      ��   �    p �       C          �    p �       C          �    p �       C          �    p �   ��fvl���H      C       �   �    � �                                                        ` � �     w       �        � � �     w          e    p �    	   w          �    p �       w          Z    p �       w          �    p �    	   w          �    p �       w      ��   �    p �       w          �    p �       w          �    p �       w          �    � �       w          �    p �       w       �   �    � �       w          �    p �   ��|R/TI
޹M.      w          �    p �       w       0        � � �                     ` � �    �      �   /     �                                                                                  ` � �                       ` � �                                  B    �                �     �         �        �                        	 H U      �   /                                        U      �   /                                           �,�*����1@2	$  �      �   /                                          �      �   /     �                                                             	               �    ` � �             0        � � �   �      �   /                                          U      �   / f                                         �      �  �                                                       �    � �    	              �    p �                  �    p �   ���÷	ۤ7/               d   �    � �     �      �   /     �                                                              �      �   /     �                                                        ` � �                       ` � �                       ` � �                  [    p � �                 \    p � �   �      �   /     �                                    	   �               @ � �                 i    p � �              �   �    p �   ��5����X"Mz,U�                 j    p � �                 �    p � �                           H                        	 H                                                                                                                                                                                                                  �                                                                                                                              �w�e�g�U            �                                                                                                                                                                    �                                                     @                             �                          �                          �                          �                          �                          �                          �              ��(� �X���r��              �                          �                                                                                                                                             d                            e                            f                            y                            z                            {                            �                            �                           �                           �              ����Sɶ�K�;�                                          "�                           '                            �                           �                           �                          m                          u                          }                          �                     ?     �                                                                                                                 
                                           ���A��I��                                                                      �                          �                          �                                                
                                                             #                           /                           ;                           >                           F                           Z                           _                           f              �����	ͦ%1�               i                           l                           y                           |                           �                           �                     
      �                           �                           �                           �                           �                           �                           �                           �                           �                           �              �]i׼�D;ҧ)               �                           �                           �                           �                           �                           �                           �                           �                           �                                                                              3                          6                          >                          E                          H              �ø����         
     c                          m                          }                          �                          �                          �                          �                          �                          �                          �                          �                          �                          �                     1     �                                                                   ����Z�Q���                                                             	                                                       �                                                        7                          P                        @                             S                          U                          X                          [                          ^                          d                     	     h              �A�4�h*̨[�S              q                          s                        M                           \                             v                          {                          �                          �                     
     �                          �                          �                          �                          �                          �                        ]                             �              ���(,C�1}��            `                             �                     
     �                          �                          �                          �                                                                              '                          .                          6                     	     F                          O                          [                     0     h                          �              ���Po�;��#              �                          �                          �                          �                          �                          �                          �                          �                                                   l                                                                                                                                                               -              �&,ﶗ��aҼ*              2                     	     8                          A                          P                     	     T                          ]                          c                          k                          r                          �                          �                          �                          �                          �                     
     �                          �              	�#_��&����a         
     �                     
     �                          �                          �                          �                     
     �                          �                          �                          �                     /     �                     
     +                          5                          @                          H                          V                          [              
��O��'9�Qǩ              c                          k                        �                             n                     	     v                     	                          	     �                     	     �                          �                     
     �                          �                          �                     	     �                        �                             �                        �                 ��S�1�� Y              �                          �                          �                        �                             �                          �                        �                                                                            
                                                         %                                                                                  !                          "              ��*Xs��K���              $                          '                          )                          +                          -                          /                          1                          3                          5                          7                          9                          :                          <                          >                          @                          B              ��l�IO=�[�              D                          F                          H                          I                          K                          M                          O                          Q                          R                          T                          V                          W                          Y                          [                          ]                          ^              �ɷ�y/�5)%��              `                          a                          b                          d                          f                          j                          l                                                  �     p                                                �                                                           �                                                    
     d                            
              ���؜�r��<�              �                                                                                                                                           @                                                                                      S                          J                                                      P                                                                                                                       ��C�üb��h                   �                           #                           2                           
                           	                                                      �                                                                        
     n                               d                                                                                  e                                                  3              �~5z�����#�y            ��������                                                                               �                                                                                                                                                                       
                                                          3                                                                           @                        
     x              ���H��|��5                                     
     �                          �                            	                           �                                                       �                                                                                  �                                                      �                                                     L                          1                          A              �W�+��wYM�A              T                          \                          Q                          a                                                                                                                                                                      !                           �                               !                        1                           �                               1                           �          �f��u�%-�zL�                                          �                                                       �                                                                                  �                                                                                  �                                                       �                                                      �                                                                      �g�?
!���;�                                           �                                                                                  �                                                                                  �                                                
     �                          +                     #     q                            �                          8                           �                            d              �Й�{����N�             I                       #     �                          =                           �                                                                                    �                           �                                                                           #     �                           �                           �                                                #     �                                          ��	��0�E&H         
     �                           �                           �                           �                           �                           �                        �                           `                                                                                     �                                                                                  �                                                                     �G�D��@U����                                                                       �                     
     �                                                                                    
                 
     �                           �                                                        l                     
     �                          �                                                
     �                                        �>��X9�U��         
     �                          �                              x                                                       �                      *                        �                        
     �                          "                              ��                                              
     �                               �                        y                                                      "�              ��~�59���
�             ����                                                     a                           f                          B                           �                            Z                          G                     #     �                            �                           #)                     P                                "                       �  /                          �                         �  -              ��N+=׼R�Ă�                                                                                              	                           �                           �                            c                                                                                                         �                 �    �  �           �M r                       �M r             �                 �    �  �           �M r                       �M r          �4߰́9�l�     }            ����      �  �           �M r                       �M r                                        �      �         �    �               �M r                        �� #�                        ω #�                                                    T                                                      d                           
                           y                                                                   s|�z) ��AN�                                            e   	                        �   
                                                                     �   "    �                  �   #    �                                                                                                    �   (    �                  �   )    �                  �       �                  �       �               	   H               x �     	   H               x �   �����V�4y�    	   H               x �     	   H               x �     	   H               x �     	   H               x �        H       �                  H       �               	   H               x �     	   H               x �     	   H               x �     	   H               x �     	   H               x �     	   H               x �                x               	   w               x �     	   w               x �     	   w               x �   �{+�sF2���$    	   w               x �     	   w               x �     	   w               x �     	   w               x �     	   w               x �     	   w               x �                                      ;    �                     =    �                     ?    �                     6    �                           �                           #                           �                                                      	              ���J��]�          I    �                      Y    �                     5    �                     g    �                     h    �                          �                                                      \                           f                      
    �                          �                      [    �                           �                           �                     r    �                �      �  ?     �    �  !��[|�C���S�                         �                                K      @  ?                                                                                                                                                                                                 *�     4   �   �                            3                     =                  *      P                  W   �   �           k      )                    @        "�N���F�     @      !                    7           7           %           K            	      	     &      "      
      
     8           �                       ,                       .                       /                          $           $                       '      A                 r      B                 s      <                 ^      F                 |                       0  #��?��R7<B�           z                       1      E                 y                 +                 E                       2      ,                 F                       3                        4      #                    9           9      .                    I           I      H                    ~           ~      I                                     2                      N           $x�7�(�:Ӛ"  N      3      !         !     O           O      &      "         "     =           =      O      #      #     �           ;      %      $      $     <           R           B           Q           P      -      %         %     G           G      $      &         &     :           :                                   �            �                        2  �                       '      '             %��6)c�c��mZ                 (      (                            )      )                	      	      *      *     
                 
      +      +                            ,      ,                            -      -                            .      .                            /      /                            0      0                            1      1                            2      2  &��wRngW<��                              3      3                            4      4                            5      5                  6      6     +      '      7      7     >      (      8      8     ?      *      9      9     A      /      :      :     J      0      ;      ;     L      1      <      <     M      4      =      =     S      5      >      >     T      6      ?      ?     U      7      @      @     V      8  '	��/j���X]�      A      A     X      9      B      B     Y      :      C      C     Z      ;      D      D     [           \           ]           _           `           a      >      E      E     b           c           d           e           f           g           h           i           j           l           m      ?      F      F     o      @      G         G     p           p      C      H      H     t     ([D�AE8��8�   D      I      I     u      G      J         J     }           }      J      K      K     �      K      L      L     �      L      M      M     �      M      N      N     �      N      O      O     �      Q      P      P     �      R      Q      Q     �      S      R      R     �      T      S      S           U      T      T     (      V      U      U     A      W      V      V     S      X      W      W     e      Y      X  )u�1;j��ΒX      X     w      Z      Y      Y     �      [      Z      Z     �      \      [      [     �      ]      \      \     6      ^      ]      ]     �      _      ^      ^     �      `      _      _           a      `      `           b      a      a           c      b      b     #      d      c      c     �      e      d      d     �      f      e      e     #      g      f      f     �      h      g      g     �      i      h  *P��K�[�z$u      h     �      j      i      i     �      k      j      j     �      l      k      k     �      m      l      l     �      n      m      m           o      n      n           p      o      o           q      p      p           r      q      q           s      r      r     %      t      s      s     *      u      t      t     >      v      u      u     C      w      v      v     P      x      w      w     U      y      x  +Svyp;x[��      x     b      z      y      y     g      {      z      z     t      |      {      {     y      }      |      |     �      ~      }      }     �            ~      ~     �      �                 �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �  ,P��.����      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     $      �      �      �     =      �      �      �     O      �      �      �     �      �      �      �     &      �      �      �     ?      �      �  -P��"�m��[s�      �     Q      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     k      �      �      �     |      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     }      �      �      �     �      �      �      �     �      �      �      �     �      �      �  .PJ���'���8�      �     1      �      �      �     F      �      �      �     a      �      �      �     s      �      �      �     �      �      �      �     �      �      �      �     2      �      �      �     G      �      �      �     c      �      �      �     u      �      �      �     �      �      �      �     
      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �  /P�E[@�}�*���      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �           �      �      �     �      �      �      �           �      �      �     ,      �      �      �     ;      �      �      �     M      �      �      �     _      �      �      �     q      �      �      �     �      �      �      �     �      �      �      �            �      �  0S[�|kX.���Ʌ      �     )      �      �      �     B      �      �      �     T      �      �      �     f      �      �      �     x      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �           �      �      �           �      �      �           �      �      �           �      �  1P�#􂪙���      �     '      �      �      �     +      �      �      �     -      �      �      �     /      �      �      �     0      �      �      �     3      �      �      �     4      �      �      �     5      �      �      �     6      �      �      �     7      �      �      �     @      �      �      �     D      �      �      �     E      �      �      �     H      �      �      �     R      �      �      �     V      �      �  2P����L�NMR�      �     W      �      �      �     X      �      �      �     Y      �      �      �     [      �      �      �     d      �      �      �     h      �      �      �     i      �      �      �     v      �      �      �     z      �      �      �     {      �      �      �     ~      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �      �     �      �      �  3P��3�,G���A      �     �      �      �      �     �      �      �      �           �      �      �     Z      �      �      �     j      �      �      �     �            �      �  �   2   3   *   +   ,   -   .   0   /   W   �   �  �  �  �  �  �  �  �  �  �  �  �  k  @  7  �  �  �  %  K  &  8  �  �  �  �  �  ,  .    	    /  $  '  r  s  ^     !  "  .  |  0  9  :  <  z  1  y    J  K  L  N  E  2  ]  ^  `  F  3  n  o  p  r  4!�㩼w���ji�  4  �  �  �  �  9  �  �  �  �  �  I  ~    N  O  =  �  �  �  �  �  ;  <  �  �  �  R  B  Q  P  G  :        �   �  �   �   �  �  �  �  �  �  �                                  !   "   #   $   %   &   '   (   7   6   ?   @   A   V   4   5   Q   8   9   :   ;   <   =   >   B   C   D   E   F   G   H   I   J   K   L   M   N   O   P   1   R   U   T   S  �  �  �  �  �              	  
                                5@m��(�v�X	                 +  >  ?  A  J  L  M  S  T  U  V  X  Y  Z  [  \  ]  _  `  a  b  c  d  e  f  g  h  i  j  l  m  o  p  t  u  }  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �    (  A  S  e  w  �  �  �  6  �  �        #  �  �  #  �  �  �  �  �  �  �            %  *  >  C  P  U  b  g  t  y  �  �  6��A| 5��  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  $  =  O  �  &  ?  Q  �  �  �  �  �  �  k  |  �  �  �  }  �  �  �  1  F  a  s  �  �  2  G  c  u  �  
  �  �  �  �  �  �  �  �  �    �    ,  ;  M  _  q  �  �     )  B  T  f  x  �  �  �  �  �  �  �          '  +  -  /  0  3  4  5  6  7  @  D  E  H  R  V  W  X  Y  [  d  h  i  v  z  {  ~  �  �  �  �  �  �  �    Z  j  �  7�����O F��B   �              �      2                                                                                    
	                  �     �      �                  	                        !      1                                          #                                          
                        �      d�           �     �      P        �   ����    ll���%���������%nn%aɕ��@�@�@�%aٖ��@�@�@�%LL%�������%����������  8�� L]�ڪ��&@�����@�@%����%������%nn%@�%a㨗�@aׁ���%LL%�@�@���%������%������%���������%��%��%������%nn%LL%������%nn%aم�������@�@�@�%aׁ����@�@�@�%a㨗�@aׁ��%LL%M]}%M]}%M]}%]}%?������%nn%@@aי��Ⅳ@�@a���@aㅧ�@�%@@aƖ��@LL@a��@�@�@�@nn%LL%�@�@���%������%nn%aŕ������@a払����ŕ������%aՁ��@a��%a⤂����@a㨗��%a㨗�@aƖ��%LL%�@�@���%������%nn%aׁ���@�@�@�%a㨗�@aÁ�����%LL%�@�@���%������%nn%aי������@M�������@��K�@M����@���Ö���k@����]]%LL%�@�@���%lBFw�%lBFw�l���`�K�%@@aƖ��@LL@a��@�@�@�@nn@@aי��Ⅳ@�@a���@aㅧ�@�  9�4;x �X���O@z@@�@�@�@��@�@���@�@�@�����@�@LLM]}\����\������\���\������\���������\������������\������������\�����������\����������\������]}a��Ɩ��@aaÖ������@aÖ���@aÙ������ā��@M�zaŕ������@a払����ŕ������a��@aɕ��@�@�@�a҉��@�aӅ����@aԅ����@�@�@�@aՁ��@a��aׁ���@�@�@�aׁ����@�@�@�aי������@M�������@��K�@M����@���Ö���k@����]]aم�������@�@�@�aٖ��@�@�@�a≩�@a⤂����@a㨗��a㉣��@Ma㨗�@aÁ�����a㨗�@aƖ��a㨗�@aׁ��a㨗�@aׁ���ll���l���`�K�mm�����m������nn�����M]@������K@������������������������M]@������K@  :"�*Y��̃�c����������������������������������������M]@������K@�����������M]@������K@�����������Ó���Ƣ���Ö�����Ù���Ƣ���Ù���Ƣ���������������������������������������ř���@���������ǉ������@Ö���������@����@`@����������|�����K��������������������������������������@@@��������������������������M]�����������������������������������������������������������������������������������������������������@����������@�����@�@�@�@����@�@�@�@�@�@����@�@����@�@����@�@������������@BFw� /?/O_o�/O%O%oo&O??_7  ;�I$̎�&}/aӃ?OD��_PY_oO�����`��/�   	�      �      �      �   ���������������������������������\����@@@\�����@@\����@@@\����@@@\���@@@@\����@@@\����@@@@@@@@@@@��������                                                                                                                ��������@@��\����@@@@@            @@@@@@@@@@  � ����     @      �               ���������@�������������@  ���Ka��������@@    @           @       @      @  @                                                                        <��@{�n��o                                                                                                                                                                                                                       \�@@@@@@@@                   �������@@@@@@@@@@@@@@@@@@@@@@@\����@@@@@@@@@@@@@@@@@@@@@@@@@��������@@@@@@@@@@@@@@@@@@@@@@\����@@@@@@@@@@@@@@@@@@@@@@@@@��������@@@@@@@@@@@@@@@@@@@@@@\����@@@@@@@@@@@@@@@@@@@@@@@@@��������@@@@@@@@@@@@@@@@@@@@@@\����@@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@�����@@@@@�����  =�6�`������@@@@@������@@@@�������@@@m������@@@mm�����@@@��������@@���������@���������@���������@���������@���������@��������������������������������������������������������������������������������                �����������������@        �������������������������   
�             �   ���������@�������������������@�����������������������������@�������@@@���������@�������������������������������������������������@�������������������������������������������������������������@����������     
`            �        >�t@"(�y���      K            �       ���������@�����������������@@@@@@@@���������@�����������������@@@@@@@@���������@�����������������@@@@@@@@���������������������������@@@@@@@@�����������\����@@@\����@@@@@@@@@@@���������������@@@@@@@@@@@@@@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��������@@@@@@@@@@@@@@@@@@@@@@          P      @@       �        �����  ������������    �@@@@@@@@@@@@@�@@@@��������@@����������\����@@@\����@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ?�W�������KQ@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�����������������������������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����������������������@@@@�������@@@��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@    ���    ��<    �� @ ��                                                                 �H             f  v   j  �   j  �   j  �     �     �                 %   .    @v`f[_���&j�      c                                            �     �                             �   #  �            n   �   l����         �   #  �   o         o         o         o         o         n   �   l����       o         !  �        q                  #  �            a                #  �           �     �         	     !   #  �            	        �   q             3         !         3                
     "   #  �     A�<�@��D��0~         
        !   #  �                             �         o                     n   �   l����         �   #  �   n   �   l����       o                 i          V   	   =   	                         o                     n   �   l����       o                �               *  f            #   >   q           $     %   a         
                o               n   �   l����                      n   �   l����       o     Ba�!7��I��b	              i          V   	   =   	             �            o                     n   �   l����       o           �           *  f                o               n   �   l����                      n   �   l����         �   #  �   n   �   l����       o           �           *  f                o               n   �   l����         �   #  �                     n   �   l����         �   #  �   n   �   l����         �   #  �   n   �   l  C/MVâϯ�s�<����       o         !  �        q                  #  �        &   a                #  �           �     �              !   #  �                    �   q             3         !         3                     "   #  �                    !   #  �                             �         o                     n   �   l����       o           '   N      K      K      #  [         o               n   �   l����       o        DT��o}��s ��     (   N      K      K      #  X         o               n   �   l����       o           )   N      K      K      #  b         o               n   �   l����       o           )   N      K      K      #  �         o               n   �   l����       o           *   N      K      K      #  +         o               n   �   l����       o           +   N      K      K      #  J         o               n   �   l����       o           +   N  E�/�n�ݿ��Z�      K      K      #  �         o               n   �   l����                      n   �   l����       o         !  �        q                  #  �        ,   a                #  �           �     �              !   #  �                    �   q             3         !         3                     "   #  �                    !   #  �                             �         o                     n   �   l����       o  F8w��Ȫv��S"           '   N      K      K      #  [         o               n   �   l����       o           (   N      K      K      #  X         o               n   �   l����       o           -   N      K      K      #  b         o               n   �   l����       o           .   N      K      K      #  �         o               n   �   l����       o           /   N      K      K      #  +         o               n   �   l����       o           G�5&y���\�:  0   N      K      K      #  J         o               n   �   l����       o           1   N      K      K      #  �         o               n   �   l����                      n   �   l����       o                 f            �            o                     n   �   l����       o           (   N      K      K      #  [         o               n   �   l����       o           '   N      K      K      #  X         o               n  H����wt�2�Y   �   l����       o           2   N      K      K      #  b         o               n   �   l����       o           3   N      K      K      #  �         o               n   �   l����       o           /   N      K      K      #  +         o               n   �   l����       o           4   N      K      K      #  J         o               n   �   l����       o           4   N      K      K      #  �         o               n   �   l����  I"��Q��
��                      n   �   l����       o                 f            �            o                     n   �   l����       o           (   N      K      K      #  [         o               n   �   l����       o           '   N      K      K      #  X         o               n   �   l����       o           -   N      K      K      #  b         o               n   �   l����       o           3   N      K      K      #  �         o  J^=�ᓣ���Z�%               n   �   l����       o           5   N      K      K      #  +         o               n   �   l����       o           6   N      K      K      #  J         o               n   �   l����       o           2   N      K      K      #  �         o               n   �   l����                      n   �   l����       o         !  �        q                  #  �        7   a                #  �           �     �           K����俌qR,     !   #  �                    �   q             3         !         3                     "   #  �                     !   #  �                              �         o                  !   n   �   l����       o                 g       	   =              =              W      K      K      #  [         o               n   �   l����       o                 e       	   =              =              W      K      K      #  X        LN���d34���   o               n   �   l����       o                 h       
   =              =              W      K      K      #  b         o               n   �   l����       o                 m       
   =              =              W      K      K      #  �         o               n      l����       o           
      ]       	   =                r            o                  "   n     l����       o                 i          V   	   =         MLG׹�$�
)x�M       W      K      K      #  +         o               n     l����          #      "      n     l����         �   #  �   n     l����       o           
      ]       	   =              =              W      K      K      #  +         o                  #      n     l����         �   #  �   n     l����       o                 `          =              =              W      K      K      #  J         o               n     l����       o     N�)I��]�              l          =              =              W      K      K      #  �         o                  !      n     l����         �   #  �            n  	   l����       o                 c            �            o                  $   n  
   l����       o                 e       	   =              =              W      K      K      #  [         o               n     l����       o                 g       	   =              =     OJq"����t�           W      K      K      #  X         o                  $      n     l����         �   #  �                  n     l����         �   #  �      %   o         o                  !  �     �   >   �  �           L      N        �   a          
          !  �     �   >   �  �           L      N        �   a          
          !  �     �   >   �  �           L      N        �   a          
          !   /   %  �              P����!ϋ# �7   %  �   n           %  �   P           %  �                                 %         e  v   f  -   j  �   j  �   j  �   g  k     �     �                 %   .        c                                            �     �                             �   #  �            n     l����         �   #  �   o         o         o         o         o         n     l����       o         !  k   #  �     9   #  �              QY���q`M�        �     :   	      	     �       3                     	     �     �   >   #  �     �     �   4   #  �            	        �     :              �     �     �   4   >   #  �      
        �     :   	           �       3                          �     �   ?   #  �     �     �   4   #  �      
                             �   q         !  �      !  �   q   �           �   #  �     �   L      a                  R��=�x�O���2  �   >   q   �           ;        �   /   #  �   L      a                   p  �   !  @   q   )         #  �   !  �   q   �              <     �              <   #  �                    �   #  �                    �   #  �     �   L      a                     �     �   >   q   )        <     �   4   L        $      a         
          p  �         o               n      l����       o         !  @     ;   N      K      K  S�[���҇��s        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  W             K               *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7  T�X�:���_R%        %   *   
                     K      K      #  ?         o               n  #   l����       o           ?   K      K        ?   K               o                     n  $   l����       o           ?   K      K      K        �      ,   `         K      *   3            �   %   -   p        �   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �  UT��<��ǻ�      �  �           L      N        �   a          
          c  )             K               *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                       ?   K               o                     n  %   l����       o           �      ,   `         K      *   3            �   %   -   p        �   %  �          !  �     VN����������  �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  C                 �          #  �            *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                     !  �   !  �   q   �         !  �   q   �        W&����I�S�h     @   a                  A   >   q   �           B   a                   !  �   q             3          #  7   p  �         o                        n  &   l����         �   #  �   n  '   l����       o         !  @     �      ,   `         K      *   3            �   %   -   p        �   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �     X8�P$���6�M�        L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                     V   	     r            o                     n  (   l����       o           �      ,   `         K      *   3            �   %   -   p        �   %  �          !  �     �      %  �        Y
����/K�2�r   %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  C                 �          #  �            *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                     !  �   !  �   q   �         !  �   q   �           C   a           Z�g/�N*+�Z��         D   >   q   �           B   a                   !  �   q             3          #  7   p  �         o                        n  )   l����         �   #  �            n  *   l����         �   #  �   n  -   l����       o         !  w   !  7   q   !               #  �        E   a                #  �           �     �              "   #  �                    �   q             3         !         3                     "  [G?b�\aP��
�   #  �                    !   #  �                             �         o                      n  .   l����       o         !  �     �               *  �            F   >   q   �        $     G   a         
          !  �   !  �     �               *  �               >   q   �        $     H   a         
          !  �   !  �     w               *  �            �   >   q   �        $     I   a         
          !  �  \�� ��������   !  7   q   !        �      ,   `         K      *   3            �   %   -   p           %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  w                      *   
      %   *            ,   `          �            �         !     �   #   7     >   %   *   
         "      !        �  ]�^�>g�gslֱ   #   7        %   *   
         "            p  �   p  �   p  �         o                         n  /   l����         �   #  �   n  2   l����       o         !  @     T   K      K        V   K      K      /     U   K      K      /     S   K      K      /   K      K        u   K      K        t   K      K      /   M      L      L        J   L      L        �      ,   `         K      *   3            �   %   -   p           %  �      ^%s��}��,ygx      !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  W             K               *   
      %   *            ,   `          �            �         #     �   #   7     >   %   *   
         $      #        �   #   7        %   *   
         $            K      K      #  ?         o               n  _7���J��aB3�  5   l����       o           ?   K      K        ?   K               o                  %   n  6   l����       o           �      ,   `         K      *   3            �   %   -   p        �   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  C                 �          #  �            *  `�٦�>"�7���   
      %   *            ,   `          �            �         &     �   #   7     >   %   *   
         '      &        �   #   7        %   *   
         '            !  �   !  �   q   �         !  �   q   �           K   a                  L   >   q   �           B   a                   !  �   q             3          #  7   p  �         o                  %      n  7   l����         �   #  �   n  :   l����       o         !  w   !  a�Tn�� �\T��  7   q   !               #  �        E   a                #  �           �     �         )     "   #  �      (      )        �   q             3         !         3                *     "   #  �      +      *        !   #  �      +         (              �         o                  ,   n  ;   l����       o         !  �     �               *  �            F   >   q   �        $     G   a         
          !  �   !  �     bO��d��.1A�  �               *  �               >   q   �        $     H   a         
          !  �   !  �     w               *  �            �   >   q   �        $     I   a         
          !  �   !  7   q   !        �      ,   `         K      *   3            �   %   -   p           %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �          c��u��L1�g��   L      N        �   a          
          c  w                      *   
      %   *            ,   `          �            �         -     �   #   7     >   %   *   
         .      -        �   #   7        %   *   
         .            p  �   p  �   p  �         o                  ,      n  <   l����         �   #  �                  n  @   l����         �   #  �      /   o         o                  !  �     �   >   �  �     d݅l*�F]X�qDS        L      N        �   a          
          !  �     �   >   �  �           L      N        �   a          
          !  �     �   >   �  �           L      N        �   a          
          !   /   %  �            8   %  �   n           %  �   P           %  �         !   /   %  �          !  @   q   )        M   L      N            a          
          !  7   q   !        M   L      N           a          
               e�B~�֐X�æV&                     /         e  -   f  �   j  �   j  �   j  �   g  %   g  K     �     �                 %   .        c                                            �     �                             �   #  �            n  E   l����         �   #  �   o         o         o         o         o         n  V   l����       o         !  %   !  }     K   K      M      L      L        �      ,   `         K      *   3            fǨ���Ci��r�  �   %   -   p        �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          a  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
         	              �   #   7        %   *   
         	                  o               n  Y   l����       o     gm2�_���y/�k        ?   K      K      K      !  %     K   K      K      K        �      ,   `         K      *   3            �   %   -   p        O   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �             K               *   
      %   *            ,   `          �            �         
     h*��|������  �   #   7     >   %   *   
               
        �   #   7        %   *   
                     K      K      #  &         o               n  Z   l����       o           &   K      K        K   K      K               o                     n  [   l����       o           �      ,   `         K      *   3            �   %   -   p        �   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L     i!�Ѭ���O�   N        �   a          
          "  �      �  �           L      N        �   a          
          c  C                 �          #  �            *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                     !  �   !  �   q   �         !  �   q   �           @   a                  A   >   q   �           B   a           j��k���M�Ti          !  �   q             3          #  8   p  �         o                        n  \   l����         �   #  �   n  _   l����       o           �   L      N      K        &   K      K      /   M      L      L      #  �         o                              n  c   l����         �   #  �         o         o                  !  �     �   >   �  �           L      N        �   a          
          !  �     �   >   �  �        k�;��ğX���g     L      N        �   a          
          !  �     �   >   �  �           L      N        �   a          
          !   /   %  �            N   %  �   n           %  �   P           %  �         !   /   %  �               #  &   !  8   q   "        M   L      N           a          
                                           e  �   f  �   j  �   j  �   j  �   g  �     �     �                 %   .        c             lج��F@�?&C%J                                 �     �                             �   #  �            n  h   l����         �   #  �   o         o         o         o         o         n  r   l����       o         !  �     q               *  �            R   >   q   �        $     S   a         
            �     3   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �     m�e�P��~��rt   %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
         	              �   #   7        %   *   
         	                  o               n  s   l����       o         !  �     o           n�{j����QƉ      *  �            T   >   q   �        $     U   a         
            �     V   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `     o��^���I�       �            �         
     �   #   7     >   %   *   
               
        �   #   7        %   *   
                           o               n  v   l����       o         "  M         �   L      N      K      K      *  M                o               n  w   l����       o         !  �     n               *  �            W   >   q   �        $     X   a         
            �     Y   N      K      K        �      ,  p�]�a�f���   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
        q^��Ʊg<|6Ya                     o               n  x   l����       o         !  �     m               *  �            O   >   q   �        $     Z   a         
            �     [   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        r�Ɗ�����E�  �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                           o               n  y   l����       o         !  �   q   �      !  \   c  �              !  �   !  �      %   ?         %   @           ]   %   ?            ^   %   @            _   #   V   !   @   q         !   ?  s�9�����nd   q         !   V   q         c  �              p  �   !  �   q   �      !  `   c  �              !  �   !  �      %   ?         %   @           a   %   ?            b   %   @            _   #   V   !   @   q         !   ?   q         !   V   q         c  �              p  �   !  �   q   �      !  �   q   �         !      q   �           c   a                  d   >   q   �           I   a                   p  �                #  ,         o  t��
X��Jbl�C               n  z   l����       o         !  �   !  ,   q            !      q   �           C   a                  D   >   q   �           e   a                   !      q   �      !  �        f   >   q   �           E   a                   !      q   �      !  �        g   >   q   �           E   a                   !  �                            *  �            h   >   q   �        $     i   a         
            �     j  uz��N�+�A[��   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       vF���'��C�X�  �   #   7        %   *   
                           o               n  {   l����       o         !  �     l               *  �            k   >   q   �        $     l   a         
            �     m   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �     w��&o:�F%t	L   �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                           o               n  |   l����       o         !  �   #       9   #                           :   	                  3                               �   >   #    xk�-�X+�g �^          �   4   #                           :                        �   4   >   #                     :   	                  3                               �   ?   #            �   4   #                                        !  �      q            !      q   �           Y   #       Y   L      a                  Y   >   q   �                   Y   /   #     L      a                   !      q  y�5�vd���M~   �      !  �           >   q   �           ;           /   #     L      a                   !      q   �      !  �           >   q   �           ;           /   #     L      a                   !  .   q            #     !      q   �           #          L      a                             >   q           n        4   L        $      a         
          p           o               n  }   l����       o         !  zԍNK��J��  �   q   �         #     !  .   q           n   #          L      a                             >   q   �        o        4   L        $      a         
            �   !  .   #       n   #                  :                        �   4   >   #                     :   	                  3                               �   ?   #            �   4   #                                             {��*���R�     N      p     K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                    |�m��$�'�h>I     �   #   7        %   *   
                           o               n  ~   l����       o         !  �     k               *  �            O   >   q   �        $     Z   a         
            �     [   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �  }?M��7�E�w���      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                           o               n     l����       o         !  �     j               *  �            F   >   q   �        $     p   a         
            �     -   N      K      K  ~���HG��::��        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �               �   #   7     >   %   *   
         !               �   #   7       ��ʷh[�q�[A   %   *   
         !                  o               n  �   l����       o         "  M         �   >     �   L      N      K      K      *  M                o               n  �   l����       o         !  �     i               *  �            W   >   q   �        $     X   a         
            �     Y   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  � �er/ԱT(�  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         "     �   #   7     >   %   *   
         #      "        �   #   7        %   *   
         #                  o               n  �   l����       o         !  �     h              ������EX�   *  �            O   >   q   �        $     Z   a         
            �     [   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `         �9�|3WW��ӄ�   �            �         $     �   #   7     >   %   *   
         %      $        �   #   7        %   *   
         %                  o               n  �   l����       o         !  �     g               *  �            q   >   q   �        $     r   a         
            �     s   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \  �hU
S���j-�Z\      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         &     �   #   7     >   %   *   
         '      &        �   #   7        %   *   
         '                  o               n  �   l����       o         !  �     f               *  �            t  ��M�������   >   q   �        $     u   a         
            �     v   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �     ��(>q򌩭�?      (     �   #   7     >   %   *   
         )      (        �   #   7        %   *   
         )                  o               n  �   l����       o         !  �     e               *  �            O   >   q   �        $     Z   a         
            �     [   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -  ���>o�N��l��]           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         *     �   #   7     >   %   *   
         +      *        �   #   7        %   *   
         +                  o               n  �   l����       o         !  �     d               *  �            F   >   q   �        $  ��0�w<X�U��     p   a         
            �     -   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         ,     �   #   7  ���$͊��#�     >   %   *   
         -      ,        �   #   7        %   *   
         -                  o               n  �   l����       o         "  M            >     �   L      N      K      K      *  M                o               n  �   l����       o         !  �     c               *  �            W   >   q   �        $     X   a         
            �     Y   N      K      K        �      ,   `         K      *   3            �ӐN��o�F2F  �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         .     �   #   7     >   %   *   
         /      .        �   #   7        %   *   
         /                  o           ��*�%�] {Ԋ      n  �   l����       o         !  �     b               *  �            O   >   q   �        $     Z   a         
            �     [   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �     �
��w61�֔1                   *   
      %   *            ,   `          �            �         0     �   #   7     >   %   *   
         1      0        �   #   7        %   *   
         1                  o               n  �   l����       o         !  �     a               *  �            w   >   q   �        $     x   a         
            �     )   N      K      K        �      ,   `         K      *   3            �   %   -   p        �=�n����/�  =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         2     �   #   7     >   %   *   
         3      2        �   #   7        %   *   
         3                  o               n  �   l����      �����l+@G�6   o         !  �     `               *  �            y   >   q   �        $     z   a         
            �     {   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *  �[)�2?v �����   
      %   *            ,   `          �            �         4     �   #   7     >   %   *   
         5      4        �   #   7        %   *   
         5                  o               n  �   l����       o         !  �     _               *  �               >   q   �        $     |   a         
            �     2   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  ���\L��i�  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         6     �   #   7     >   %   *   
         7      6        �   #   7        %   *   
         7                  o               n  �   l����       o         !  �     �}�&����&D�     q                  #          }   a                #                  �         9     !   #        8      9           q             3         !         3                :     "   #        ;      :        !   #        ;         8                       o                  <   n  �   l����       o         !  A     �               *  A            F   >   q   *        $     ~   a         
                o        �^���Cd��B         n  �   l����          =      <      n  �   l����         �   #  �   n  �   l����       o         !  A   q   *         #          q           4   #          L      a                         o                  =      n  �   l����         �   #  �   n  �   l����       o         !  A   #       4   #              >             :   	      ?            3                     ?          �   >   #            �   4   #    �	d|����k��
      >      ?             :         B               �   4   >   #        @             :   	      A            3                     A          �   ?   #            �   4   #        @      A         B                 !  �      q   *         !      q   �           .   #       .   L      a                  .   >   q   �                   .   /   #     L      a                   !      q   �      !  �          ���D�Ն���t�   >   q   �           ;           /   #     L      a                   !  .   q            #     !      q   �           #          L      a                             >   q           n        4   L        $      a         
          p           o               n  �   l����       o         !  �   q   �         #     !  .   q           n   #          L      a                             >   q   �        o       ��!o�����m�   4   L        $      a         
            �   !  .   #       n   #                  :         E               �   4   >   #        C             :   	      D            3                     D          �   ?   #            �   4   #        C      D         E                         N      p     K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  ��G	l�m+�C=��  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         F     �   #   7     >   %   *   
         G      F        �   #   7        %   *   
         G                  o               n  �   l����       o         !  �     ^              ����̲��EZ��   *  �               >   q   �        $     �   a         
            �     �   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `         �9�|3WW���   �            �         H     �   #   7     >   %   *   
         I      H        �   #   7        %   *   
         I                  o               n  �   l����       o         !  �     ]               *  �            O   >   q   �        $     Z   a         
            �     [   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \  �hU&S҈�ju�A�      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         J     �   #   7     >   %   *   
         K      J        �   #   7        %   *   
         K                  o               n  �   l����       o         !  �     \               *  �            F  ��MX{���u^   >   q   �        $     p   a         
            �     -   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �     ��(>p����?      L     �   #   7     >   %   *   
         M      L        �   #   7        %   *   
         M                  o               n  �   l����       o         "  M         �   >     �   L      N      K      K      *  M                o               n  �   l����       o         !  �     [               *  �            W   >   q   �        $     X   a         
            �     Y   N      K      K        �      ,   `         K  ����7~��      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         N     �   #   7     >   %   *   
         O      N        �   #   7        %   *   
         O           �>I�� n�,����         o               n  �   l����       o         !  �     Z               *  �            O   >   q   �        $     Z   a         
            �     [   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a         ����7�����O1   
          c  �                      *   
      %   *            ,   `          �            �         P     �   #   7     >   %   *   
         Q      P        �   #   7        %   *   
         Q                  o               n  �   l����       o         !  �     Y               *  �            �   >   q   �        $     �   a         
            �     �   N      K      K        �      ,   `         K      *   3            ��aKC�[L���2&  �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         R     �   #   7     >   %   *   
         S      R        �   #   7        %   *   
         S                  o           ���J���_`~t�      n  �   l����       o         !  �     X               *  �            �   >   q   �        $     �   a         
            �     �   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �     �
�aal��941                   *   
      %   *            ,   `          �            �         T     �   #   7     >   %   *   
         U      T        �   #   7        %   *   
         U                  o               n  �   l����       o         !  �     W               *  �            O   >   q   �        $     Z   a         
            �     [   N      K      K        �      ,   `         K      *   3            �   %   -   p        �=���vʲ	5�`  =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         V     �   #   7     >   %   *   
         W      V        �   #   7        %   *   
         W                  o               n  �   l����      �����lD Jö   o         !  �     V               *  �            F   >   q   �        $     p   a         
            �     -   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  �                      *  �[)�v ��1ĥ   
      %   *            ,   `          �            �         X     �   #   7     >   %   *   
         Y      X        �   #   7        %   *   
         Y                  o                              n  �   l����         �   #  �      Z   o         o                  !  �     �   >   �  �           L      N        �   a          
          !  �     �   >   �  �           L      N        �   a          
          !  �     ����`�aou"�  �   >   �  �           L      N        �   a          
          !   /   %  �            P   %  �   n        Q   %  �          !  �   %  �            #   %  �   P           %  �         !   /   %  �          !  ,   q           M   L      N           a          
          !  .   q           M   L      N           a          
                                  Z         e  �   f  �   j  �   j  �   j  �     �     �              �;�K鵠��z�U     %   .        c                                                 �                             �   #              n  �   l����         �   #  �   o         o         o         o         o         n  �   l����                !  �   %   /   �        �   %  �  �      !   R   q              L      N        �   a          
            �   %  �   L        �   %  �   
         �   %  �  �        �  �        �         
     ��������E�~  �   %  �   
        �      #   7   %   /   �         /   �        �   	           �          %   *   �        �  �      %   *   �        �   
       %   *   �         �   L      %   *  c                        
           %  
               %  
         !  
   q   �      c                  
         %  �   �        �   %  �   �        �   %   /   �        s   #  #   j     l����       !   /   c                k     l����          /  �+63J4W����	   �      #   7      /   �        �   
                     /   �      #   7   !  	      /   �      c                   	               	               n  �   l����       o           #                    o                     n  �   l����       o           �      ,   `         K      *   3            �   %   -   p        �   %  �          !  �     �      %           %   -   \      "   -   f   �   -           L      N        �   a  �W)|��9�x�f          
          "        �             L      N        �   a          
          c  x             K               *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                     K      K      #  $         o               n  �   l����       o                  !  �   %   /   �        s   #  #     �   %  �  �      !   R   q  ����"V` U_b�              L      N        �   a          
            �   %  �   L        �   %  �   
         �  �        �              �   %  �   
        �      #   7   %   /   �         /   �        �   	           �          %   *   �        �  �      %   *   �        �   
       %   *   �         �   L      %   *  c                                �   %   /   �        �   #   �     �   %   .        c                     /   �      #   7  �F�;3�0�Τ�      /   �        �   
                     /   �      #   7   !  	      /   �      c                                 �  �        �                 #  #                    �   %   -   D        E   #   �     �   %   .        c                    �   �        �   *   2       !     �   `   "   #   �     %   #   �     �   %   .        c                                 o                        n  �   l����       o           #     ���1"򑔶�%x                 o                     n  �   l����       o         !       �               *              �   >   q   �        $     �   a         
                 ;   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %           %   -   \      "   -   f   �   -           L      N        �   a          
          "        �             L      N     �L&����zn��     �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                           o               n  �   l����       o         !  ^   q   <         #     !  L   q   0        5   #          L      a                             >   q   <        �        4   L        $      a     �C/�_9��q���      
                o               n  �   l����       o         !     #        !      !  '   #                "             ;   N      K      K      *  '                                 '          K      K        �   K      	                                !     #        !      #                 '          K           /   K      K      *  '                                o               n  �   l����       o        ��P�����p     :   N      K      K      #  r         o               n  �   l����       o           ;   N      K      K      #  s         o               n  �   l����          $      %      n  �   l����       o           s   K      K        !   K               o                  &      '      &         $      n  �   l����       o           '   K      K      #     !  �           #                  [   N            (          "   
     ��Z69�P�pn3�   )      (        �   !  	      c                   )                 4     "   K                  /   #                  [   N            *          !   
      +      *        �   !  	      c                   +            M      #     >     r   K      K        "   K      /   #     !  ^           #                  �   N            ,          "   
      -      ,        �   !  	      c                   -     �!�@�>|tHf�              4   M           �      4   #     >         q   <        �        L           L        �     �   c                K         #                  !   
      .     �   !  	      c                   .            K      K      K      #  s         o               n  �   l����       o           s   K      K        !   K      	         o                  /   n  �   l����       o           r   K      K        s   K  �	�C	��4�J9>*      K      /   K      K      #  r         o               n  �   l����       o           !   K      #       r   K      K      #     !  ^   q   <      #     !  �   #                  �     �   /   N            0          !   
      1      0        �   !  	      c                   1                         �   N            2          !   
      3      2        �   !  	      c                   3                   �+ָ�gD��X�J     4   #       :   #     !     q   �           q   <           M      L      a                     M              /   #     >     ;      q   �                    L      a                           /   #     >   #          M           M      /   N      #             �   N                 4     �   N           4   M           q   �                M      >   q   <               L      a                     ���"%�oV�@>KU     /   #        4                 #     !     !  ^   q   <               #        q   �              �              5     �   #        6      5           #        6                 #          L      a                             >   q   <        �        4   L        $      a         
          p           o               n  �   l����       o           r   K      K        "   K      /   K      K      #  r  ���0�T����S         o                  /      n  �   l����         �   #  �   n  �   l����          %      '      n  �   l����         �   #  �   n  �   l����                      n  �   l����       n  �   l����       o         !  ^   #       �   #                  :         9               �   4   >   #        7             :   	      8            3                     8          �   ?   #            �   4   #        7      8     �esR2GT��o      9                 !     q   �               #        q   <           #          L      a                             >   q   �        o        4   L        $      a         
               p     !  ^   #       �   #                  :         <               �   4   >   #        :             :   	      ;            3                     ;          �   ?   #            �   4   #        :     �p��<�]���d   ;         <                         N      p     K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %           %   -   \      "   -   f   �   -           L      N        �   a          
          "        �             L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         =     �   #   7  �㸺.��îc     >   %   *   
         >      =        �   #   7        %   *   
         >                  o               n  �   l����       o         !       T               *              O   >   q   �        $     Z   a         
                 [   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %           %   -   \      "   -   f   �   -           L      N  ��2�0�-Ċ        �   a          
          "        �             L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         ?     �   #   7     >   %   *   
         @      ?        �   #   7        %   *   
         @                  o               n  �   l����       o            A      !  �   %   /   �        s   #  #     �   %  �  �      !   R   q             �jd@ʩe�b�   L      N        �   a          
            �   %  �   L        �   %  �   
         �  �        �         C     �   %  �   
        �      #   7   %   /   �         /   �        �   	      D     �          %   *   �        �  �      %   *   �        �   
       %   *   �         �   L      %   *  c         D         E      C        �   %   /   �        �   #   �     �   %   .        c                     /   �      #   7      /   �     ��y�m�Bc���M     �   
      F      E         /   �      #   7   !  	      /   �      c                   B      F        �  �        �         G        #  #      B      G        �   %   -   D        E   #   �     �   %   .        c                    �   �        �   *   2       !     �   `   "   #   �     %   #   �     �   %   .        c                     B            o               n  �   l����       o           #                    o     �Jr�))�e��               H   n  �   l����         �   #  �   n  �   l����       o           >     �            o                  I   n  �   l����       o         !  $   q           �      ,   `         K      *   3            �   %   -   p        �   %  �          !  �     �      %           %   -   \      "   -   f   �   -           L      N        �   a          
          "        �             L      N        �   a          
          c  ���R��qc�o�  5                      *   
      %   *            ,   `          �            �         J     �   #   7     >   %   *   
         K      J        �   #   7        %   *   
         K                  o               n  �   l����       o           �      ,   `         K      *   3            �   %   -   p        �   %  �          !  �     �      %           %   -   \      "   -   f   �   -           L      N        �   a          
  �Ͽ���יm���#          "        �             L      N        �   a          
          c  x             K               *   
      %   *            ,   `          �            �         L     �   #   7     >   %   *   
         M      L        �   #   7        %   *   
         M            K      K      #  $         o               n  �   l����          N      I      n  �   l����       o           >     �            o                  O   n  ����n��s1����  �   l����       o         !       S               *         #        >   q   �        $     �   a         
                 �   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %           %   -   \      "   -   f   �   -           L      N        �   a          
          "        �             L      N        �   a          
          c  �            �q�Zukr��yyD�            *   
      %   *            ,   `          �            �         P     �   #   7     >   %   *   
         Q      P        �   #   7        %   *   
         Q                  o               n  �   l����          N      O      n  �   l����       o           >     �            o                  R   n  �   l����       o         !       R               *         #        >   q   �        $     �   a         
         �09T� �J�C�          �   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %           %   -   \      "   -   f   �   -           L      N        �   a          
          "        �             L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         S     �   #   7     >   %   *   
         T  �1Ԓ�M:J�i      S        �   #   7        %   *   
         T                  o               n  �   l����       o         !       Q               *         #        >   q   �        $     �   a         
                 �   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %           %   -   \      "   -   f   �   -           L      N        �   a          
      �2������N      "        �             L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         U     �   #   7     >   %   *   
         V      U        �   #   7        %   *   
         V                  o                  R      n  �   l����         �   #  �      N         H      n  �   l����         �   #  �   n  �   l����                      n  �   l����      ���gv_����     �   #  �   n  �   l����       o         !  $   q           �      ,   `         K      *   3            �   %   -   p        �   %  �          !  �     �      %           %   -   \      "   -   f   �   -           L      N        �   a          
          "        �             L      N        �   a          
          c  5                      *   
      %   *            ,   `          �            �         W     �   #   7     �<��5�-f�ֽ�  >   %   *   
         X      W        �   #   7        %   *   
         X                  o               n  �   l����                      n  �   l����         �   #  �   n  �   l����          Y      !  �   %   /   �        �   %  �  �      !   R   q              L      N        �   a          
            �   %  �   L        �   %  �   
         �   %   /   �      j     l����       !   /     �        #  #   c                k    Ņ��@t��   l����       !  �      %  �   0      %  �   @         /   �      #   7      /   �        �   
      [      /   �      #   7   !  	      /   �      c                   Z      [         Z                     n  �   l����         �   #  �      \   o         o                  !  	     �   >   �  	           L      N        �   a          
          !  	     �   >   �  	           L      N        �   a          
          !  	     �   >  ƓAK�G�$�A"�   �  	           L      N        �   a          
          !   /   %  	            �   %  	   n           %  	   P           %  	         !   /   %            !  /   q           M   L      N           a          
               #  $     �   #  '     �   #  r     �   #  s   !  ^   q   <        M   L      N           a          
                                  \         e  �   f  x   j  �   j  �   j  �     �     �        ���-w
��Kr�W�           %   .        c                                                  �                             �   #               n  �   l����         �   #  �   o         o         o         o         o         n  �   l����       o           �   K      K        "   K      /   K      K      #  �         o               n  �   l����       o         "  M         �   K      #  #           #     �   L      N      	           #     ț�����~a4�  �   K      	      	              �   L      N      #  #      	              #   M      L        �   4     �   �   N      A        �   L      N      K      K      *  M                o               n  �   l����       o           Y   K      K        "   K      /   K      K      #  Y         o               n  �   l����       o         "  Z         Y   K      #  #           #     �   L      N      	      
     #     �   K      	  �xS�����/g�            
        �   L      N      #  #                    #   M      L        �   4     �   �   N      A        �   K      K      K      *  Z                o               n  �   l����       o           �   K      V      U         %  $       $         !  &     �   >   q   �      !  $   q   �            a                #  '     �   #  (              (        
           '      &            s              (     �   N  ʝ�c�湌qH      /   #  (     '     �   >   #  '                    $           s   G     �              '     �   ?      #  '     �   *  &            &           s   I   %  &                          '        �      !  &   @   4   M      #  %   q   �      !  |      !  )   q   �           %   #  *     %   L      a                  %   >   q   �           V        %   /   #  *   L      a                   p  &   p  %   !  )   q   �  �}�R����'      !  �        *   >   q   �           ;        *   /   #  *   L      a                   !  0   q            #  +   !  )   q   �        *   #  %     %   L      a                     +     %   >   q           n     %   4   L        $      a         
          p  *         o               n  �   l����       o         !  ,   q   �         #  +   !  0   q           n   #  %     %   L      a                     +     %   >   q  ̴�����,����(   �        o     %   4   L        $      a         
            ,   !  0   #  +     n   #  %           %     :              +     %     �   4   >   #  -              %     :   	           -       3                          -     �   ?   #  -     %     �   4   #  %                                   +        %   N      p  %   K        �      ,   `         K      *   3            �   %   -   p        =   %  �         ������[̯��   !  �     �      %  .         %   -   \      "   -   f   �   -           L      N        �   a          
          "  .      �  .           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                           o               n  �   l����       o         !  ,  ��z�h�A��Wʵ     P               *  ,            O   >   q   �        $     Z   a         
            ,     [   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  .         %   -   \      "   -   f   �   -           L      N        �   a          
          "  .      �  .           L      N        �   a          
          c  �                      *   
      %   *     ϸ�.FmcI�hш         ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                           o               n      l����       o         !  ,     O               *  ,            w   >   q   �        $     x   a         
            ,     )   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  �x1a���R"�}�  .         %   -   \      "   -   f   �   -           L      N        �   a          
          "  .      �  .           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                           o               n     l����       o         !  ,     N              ў���qQ��c�n   *  ,            �   >   q   �        $     �   a         
            ,     �   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  .         %   -   \      "   -   f   �   -           L      N        �   a          
          "  .      �  .           L      N        �   a          
          c  �                      *   
      %   *            ,   `         �8�]|4b���/+   �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                           o               n     l����       o         !  ,     M               *  ,            �   >   q   �        $     �   a         
            ,     �   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  .         %   -   \  �hUh�r����D,      "   -   f   �   -           L      N        �   a          
          "  .      �  .           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                           o               n     l����       o           �   K      K        "   K      /   K      K  ������|&r      #  �         o               n     l����       o           �   K      V      U         %  $       $         !  &     �   >   q   �      !  $   q   �            a                #  +     �   #  (              (        
           +      &            s              (     �   N      /   #  (     +     �   >   #  +                    $           s   G     �              +     �   ?      #  +     �   *  &            ��4	������d  &           s   I   %  &                          +        �      !  &   @   4   M      #  %   !  �      q   �         !  )   q   �           2   #  *     2   L      a                  2   >   q   �           %        2   /   #  *   L      a                   !  )   q   �      !  }        *   >   q   �           �        *   /   #  *   L      a                   !  )   q   �      !  �        *   >   q   �           ;        �]0�}�z�<g�  *   /   #  *   L      a                   !  0   q            #  -   !  )   q   �        *   #  %     %   L      a                     -     %   >   q           n     %   4   L        $      a         
          p  *         o               n     l����       o         !  ,   q   �         #  -   !  0   q           n   #  %     %   L      a                     -     %   >   q   �        o     %   4   L        $      a        �*C�䓄cUV��   
            ,   !  0   #  -     n   #  %           %     :         !     -     %     �   4   >   #  /              %     :   	            /       3                           /     �   ?   #  /     %     �   4   #  %                      !              -        %   N      p  %   K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  .         %   -   \      "   -  �a�Z��8�e�ؕ   f   �   -           L      N        �   a          
          "  .      �  .           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         "     �   #   7     >   %   *   
         #      "        �   #   7        %   *   
         #                  o               n     l����       o         !  ,     L               *  ,            O   >   q   �  �A��\ɬ��r��        $     Z   a         
            ,     [   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  .         %   -   \      "   -   f   �   -           L      N        �   a          
          "  .      �  .           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         $     ڼ���<���n?h  �   #   7     >   %   *   
         %      $        �   #   7        %   *   
         %                  o               n     l����       o         !  ,     K               *  ,            F   >   q   �        $     p   a         
            ,     -   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  .         %   -   \      "   -   f   �   -          ۑ���r�et�t   L      N        �   a          
          "  .      �  .           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         &     �   #   7     >   %   *   
         '      &        �   #   7        %   *   
         '                  o               n  	   l����       o         "  M         �   K      #  #           #     �   L      N      	      (     ����$�S��r  #     �   K      	      )      (        �   L      N      #  #      )              #   M      L        �   4     �   �   N      A        �   L      N      K      K      *  M                o               n  
   l����       o           �   K      V      U         %  $       $         !  &     �   >   q   �      !  $   q   �            a                #  -     �   #  (      *        (        
      +     -      &            s  ��c
wg��7�-         +     (     �   N      /   #  (     -     �   >   #  -      *      +        $           s   G     �         ,     -     �   ?      #  -     �   *  &            &           s   I   %  &            ,              -        �      !  &   @   4   M      #  %   q   �      !  |      !  )   q   �           %   #  *     %   L      a                  %   >   q   �           V        %   /   #  *   L      a                  �|��PZ�!�?��   p  &   p  %   !  )   q   �      !  �        *   >   q   �           ;        *   /   #  *   L      a                   !  0   q            #  /   !  )   q   �        *   #  %     %   L      a                     /     %   >   q           n     %   4   L        $      a         
          p  *         o               n     l����       o         !  ,   q   �         #  /   !  0   q           n   #  %     %   L      a           ��fòm��01            /     %   >   q   �        o     %   4   L        $      a         
            ,   !  0   #  /     n   #  %           %     :         /     /     %     �   4   >   #  0      -        %     :   	      .     0       3                     .     0     �   ?   #  0     %     �   4   #  %      -      .         /              /        %   N      p  %   K        �      ,   `         K      *   3            �   %   -  �{�jkQ�̀8���   p        =   %  �          !  �     �      %  .         %   -   \      "   -   f   �   -           L      N        �   a          
          "  .      �  .           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         0     �   #   7     >   %   *   
         1      0        �   #   7        %   *   
         1                  o               n    ��GU���Aܫ   l����       o         !  ,     J               *  ,            O   >   q   �        $     Z   a         
            ,     [   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  .         %   -   \      "   -   f   �   -           L      N        �   a          
          "  .      �  .           L      N        �   a          
          c  �               �hg��J��0�Zl         *   
      %   *            ,   `          �            �         2     �   #   7     >   %   *   
         3      2        �   #   7        %   *   
         3                  o               n     l����       o           �   K      K        "   K      /   V      U         %  1       %         !  2     �   >   q   �      !  1   q   �        �   a                #  /     �   #  (      4        (     �   
      5     /      �1E��g�1f�  2            s         5     (     �   N      /   #  (     /     �   >   #  /      4      5        1           s   G     �         6     /     �   ?      #  /     �   *  2            2           s   I   %  2            6              /        �      !  2   @   4   M      #  %   !  �      q   �         !  )   q   �           Y   #  *     Y   L      a                  Y   >   q   �           %        Y   /   #  *   L     䉃��F�ά1�1t   a                   !  )   q   �      !  }        *   >   q   �           �        *   /   #  *   L      a                   !  )   q   �      !  �        *   >   q   �           ;        *   /   #  *   L      a                   !  0   q            #  0   !  )   q   �        *   #  %     %   L      a                     0     %   >   q           n     %   4   L        $      a         
          p  *         o              �J���T$a�   n     l����       o         !  ,   q   �         #  0   !  0   q           n   #  %     %   L      a                     0     %   >   q   �        o     %   4   L        $      a         
            ,   !  0   #  0     n   #  %           %     :         9     0     %     �   4   >   #  3      7        %     :   	      8     3       3                     8     3     �   ?   #  3     %     �   4   #  %      7      8     ��ٵu�2t�      9              0        %   N      p  %   K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  .         %   -   \      "   -   f   �   -           L      N        �   a          
          "  .      �  .           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         :     �   #   7     >  �V�w)�cīM7��   %   *   
         ;      :        �   #   7        %   *   
         ;                  o               n     l����       o         !  ,     I               *  ,            O   >   q   �        $     Z   a         
            ,     [   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  .         %   -   \      "   -   f   �   -           L      N        躳{�2K���/  �   a          
          "  .      �  .           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         <     �   #   7     >   %   *   
         =      <        �   #   7        %   *   
         =                  o               n     l����       o         !  ,     H               *  ,            F   >   q   �        $     p   a         
         �-s�et>`�     ,     -   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  .         %   -   \      "   -   f   �   -           L      N        �   a          
          "  .      �  .           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         >     �   #   7     >   %   *   
         ?  �1ԋ 
�:
$�5      >        �   #   7        %   *   
         ?                  o               n     l����       o           �   L      N      K      K      #  |         o               n     l����       o         !  ,     G               *  ,            O   >   q   �        $     Z   a         
            ,     [   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �     �S�"x�9��#L   %  .         %   -   \      "   -   f   �   -           L      N        �   a          
          "  .      �  .           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         @     �   #   7     >   %   *   
         A      @        �   #   7        %   *   
         A                  o               n     l����       o           b   K      V      U  �� �rL'[N�         %  $       $         !  &     �   >   q   �      !  $   q   �            a                #  0     �   #  (      B        (        
      C     0      &            s         C     (     �   N      /   #  (     0     �   >   #  0      B      C        $           s   G     �         D     0     �   ?      #  0     �   *  &            &           s   I   %  &            D              0        �      !  &   @   4  �W7{�ߨ�!A�   M      #  %   !  �      q   �         !  )   q   �           �   #  *     �   L      a                  �   >   q   �           %        �   /   #  *   L      a                   !  )   q   �      !  y        *   >   q   �           [        *   /   #  *   L      a                   !  )   q   �      !  �        *   >   q   �           ;        *   /   #  *   L      a                   !  0   q            #  3   !  )   q   �     ����K�A�~���     *   #  %     %   L      a                     3     %   >   q           n     %   4   L        $      a         
          p  *         o               n     l����       o         !  ,   q   �         #  3   !  0   q           n   #  %     %   L      a                     3     %   >   q   �        o     %   4   L        $      a         
            ,   !  0   #  3     n   #  %           %     :         G     3     �
�a*�x�3Q[
  %     �   4   >   #  4      E        %     :   	      F     4       3                     F     4     �   ?   #  4     %     �   4   #  %      E      F         G              3        %   N      p  %   K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  .         %   -   \      "   -   f   �   -           L      N        �   a          
          "  .      �  .        �ݜ�B��?b� '     L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         H     �   #   7     >   %   *   
         I      H        �   #   7        %   *   
         I                  o               n     l����       o           J   K      V      U         %  $       $         !  &     �   >   q   �      !  $   q   �            a                #  3     �   #  (     �|����A�u�}   J        (        
      K     3      &            s         K     (     �   N      /   #  (     3     �   >   #  3      J      K        $           s   G     �         L     3     �   ?      #  3     �   *  &            &           s   I   %  &            L              3        �      !  &   @   4   M      #  %   !  �      q   �         !  )   q   �           Y   #  *     Y   L      a                  Y   >   q   �  �rxT�f�؄�           %        Y   /   #  *   L      a                   !  )   q   �      !  w        *   >   q   �           ;        *   /   #  *   L      a                     X   K      K        �   K      K      4   V      U         %  1       %         !  2     �   >   q   �      !  1   q   �        �   a                #  4     �   #  (      M        (     �   
      N     4      2            s         N     (     �   N      /   #  ���D��]<!  (     4     �   >   #  4      M      N        1           s   G     �         O     4     �   ?      #  4     �   *  2            2           s   I   %  2            O              4        �      !  2   @   4   M      #  %   !  )   q   �         q   �           *   >   q   �           %        *   /   #  *   L      a                   !  )   q   �      !  z        *   >   q   �           [        *   /   #  *   L      a  ��7 �X�ό�                   !  )   q   �      !  �        *   >   q   �           ;        *   /   #  *   L      a                   !  0   q            #  5   !  )   q   �        *   #  %     %   L      a                     5     %   >   q           n     %   4   L        $      a         
          p  *         o               n     l����       o         !  ,   q   �         #  5   !  0   q           n   #  %     %   L      a        �9tR�4�Tw�               5     %   >   q   �        o     %   4   L        $      a         
            ,   !  0   #  5     n   #  %           %     :         R     5     %     �   4   >   #  6      P        %     :   	      Q     6       3                     Q     6     �   ?   #  6     %     �   4   #  %      P      Q         R              5        %   N      p  %   K        �      ,   `         K      *   3            �   %  �u' d��q�V��   -   p        =   %  �          !  �     �      %  .         %   -   \      "   -   f   �   -           L      N        �   a          
          "  .      �  .           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         S     �   #   7     >   %   *   
         T      S        �   #   7        %   *   
         T                  o               n  �{�J��.�ފ�  "   l����       o           �   K      V      U         %  $       $         !  &     �   >   q   �      !  $   q   �            a                #  5     �   #  (      U        (        
      V     5      &            s         V     (     �   N      /   #  (     5     �   >   #  5      U      V        $           s   G     �         W     5     �   ?      #  5     �   *  &            &           s   I   %  &           �A-��^��e	��   W              5        �      !  &   @   4   M      #  %   q   �      !  {      !  )   q   �           %   #  *     %   L      a                  %   >   q   �           [        %   /   #  *   L      a                   p  &   p  %   !  )   q   �      !  �        *   >   q   �           ;        *   /   #  *   L      a                   !  0   q            #  6   !  )   q   �        *   #  %     %   L      a                  ���|���I���     6     %   >   q           n     %   4   L        $      a         
          p  *         o               n  #   l����       o         !  ,   q   �         #  6   !  0   q           n   #  %     %   L      a                     6     %   >   q   �        o     %   4   L        $      a         
            ,   !  0   #  6     n   #  %           %     :         Z     6     %     �   4   >   #  7      X        %     :  �K��Tl���   	      Y     7       3                     Y     7     �   ?   #  7     %     �   4   #  %      X      Y         Z              6        %   N      p  %   K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  .         %   -   \      "   -   f   �   -           L      N        �   a          
          "  .      �  .           L      N        �   a          
          c  ���.ضuM'~�  �                      *   
      %   *            ,   `          �            �         [     �   #   7     >   %   *   
         \      [        �   #   7        %   *   
         \                  o               n  %   l����       o           |   K      K      K      h     �   #  !         o                                    n  (   l����         �   #  �     !     �         ]     �   !  "      c                   ]     ��g����bM�/�      ^   o         o                       #  !   !  "     �   >   �  "           L      N        �   a          
          !  "     �   >   �  "           L      N        �   a          
          !  "     �   >   �  "           L      N        �   a          
          !   /   %  "            �   %  "   n           %  "   P           %  "         !   /   %  .               #  |   !  0   q           M   L      N          �"�4�w�|f)   a          
                                  ^         e  x   f  5   j  �   j  �   j  �   g       �     �                 %   .        c                                            9     �                             �   #  9            n  -   l����         �   #  �   o         o         o         o         o         n  6   l����       o         !  ;     F               *  ;            O   >   q   �        $     Z  ��Q���h�.p   a         
            ;     [   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  <         %   -   \      "   -   f   �   -           L      N        �   a          
          "  <      �  <           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >  �V�w//��߻   %   *   
         	              �   #   7        %   *   
         	                  o               n  7   l����       o           �   L      N      K      K      #  y         o               n  8   l����       o         !  ;     E               *  ;               >   q   �        $     |   a         
            ;     2   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �       �,%��
Gg�      !  �     �      %  <         %   -   \      "   -   f   �   -           L      N        �   a          
          "  <      �  <           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         
     �   #   7     >   %   *   
               
        �   #   7        %   *   
                           o               n  9   l����       o         !  ��ګ�O�_O�m  ;     D               *  ;            F   >   q   �        $     p   a         
            ;     -   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  <         %   -   \      "   -   f   �   -           L      N        �   a          
          "  <      �  <           L      N        �   a          
          c  �                      *   
      %   *  ��&7��H����            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                           o               n  ;   l����       o           �   K      K        "   K      /   K      K      #  �         o               n  <   l����       o         "  M         �   K      #  #           #     �   L      N      	           #     �   K      	                    �  YD6	3z=w   L      N      #  #                    #   M      L        �   4     �   �   N      A        �   L      N      K      K      *  M                o               n  >   l����       o           �   K      V      U         %  =       $         !  ?     �   >   q   �      !  =   q   �            a                #  @     �   #  A              A        
           @      ?            s              A     �   N      /   #  A     ��n�q1�r��l   @     �   >   #  @                    =           s   G     �              @     �   ?      #  @     �   *  ?            ?           s   I   %  ?                          @        �      !  ?   @   4   M      #  >   q   �      !  |      !  B   q   �           >   #  C     >   L      a                  >   >   q   �           V        >   /   #  C   L      a                   p  ?   p  >   !  B   q   �      !  �        0�Lop�#?��  C   >   q   �           ;        C   /   #  C   L      a                   !  1   q            #  D   !  B   q   �        C   #  >     >   L      a                     D     >   >   q           n     >   4   L        $      a         
          p  C         o               n  ?   l����       o         !  ;   q   �         #  D   !  1   q           n   #  >     >   L      a                     D     >   >   q   �        o     �ͭ�ōOJ�՝�  >   4   L        $      a         
            ;   !  1   #  D     n   #  >           >     :              D     >     �   4   >   #  E              >     :   	           E       3                          E     �   ?   #  E     >     �   4   #  >                                   D        >   N      p  >   K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �     �}i�ڨ��b�   %  <         %   -   \      "   -   f   �   -           L      N        �   a          
          "  <      �  <           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                           o               n  A   l����       o           y   K      K        �v���L3 ��        z          K      K      4   V      U         %  F       %         !  G     �   >   q   �      !  F   q   �        �   a                #  D     �   #  A              A     �   
           D      G            s              A     �   N      /   #  A     D     �   >   #  D                    F           s   G     �              D     �   ?      #  D     �   *  G            G           s   I   %  G              	��lLy�x���              D        �      !  G   @   4   M      #  >   q   �      !  �      !  B   q   �           >   #  C     >   L      a                  >   >   q   �           ;        >   /   #  C   L      a                   p  G   p  >   !  1   q            #  E   !  B   q   �        C   #  >     >   L      a                     E     >   >   q           n     >   4   L        $      a         
          p  C         o           
�Ġ�8rE]��      n  B   l����       o         !  ;   q   �         #  E   !  1   q           n   #  >     >   L      a                     E     >   >   q   �        o     >   4   L        $      a         
            ;   !  1   #  E     n   #  >           >     :              E     >     �   4   >   #  H              >     :   	           H       3                          H     �   ?   #  H     >     �   4   #  >              2^8�$�F@q)�(                       E        >   N      p  >   K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  <         %   -   \      "   -   f   �   -           L      N        �   a          
          "  <      �  <           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     <�E���.���  >   %   *   
                       �   #   7        %   *   
                           o               n  D   l����       o         !  ;     C               *  ;            F   >   q   �        $     p   a         
            ;     -   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  <         %   -   \      "   -   f   �   -           L      N     錷 Ӽ�̜�2     �   a          
          "  <      �  <           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �               �   #   7     >   %   *   
         !               �   #   7        %   *   
         !                  o                              n  G   l����         �   #  �      "   o         o                  !  :     �   >   �  :          :�G(�+фa8�   L      N        �   a          
          !  :     �   >   �  :           L      N        �   a          
          !  :     �   >   �  :           L      N        �   a          
          !   /   %  :            �   %  :   n           %  :   P           %  :         !   /   %  <          !  1   q           M   L      N           a          
               #  y                           "         e  5   f  �   j  �   j  �  ]��`��)��   j  �     �     �                 %   .        c                                            J     �                             �   #  J            n  L   l����         �   #  �   o         o         o         o         o         n  U   l����       o         "  M            >     �   L      N      K      K      *  M                o               n  V   l����       o         !  M     B               *  M            W  X�55�6l%N   >   q   �        $     X   a         
            M     Y   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  N         %   -   \      "   -   f   �   -           L      N        �   a          
          "  N      �  N           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �     8(�iN��s��s           �   #   7     >   %   *   
         	              �   #   7        %   *   
         	                  o               n  W   l����       o         !  M     A               *  M            O   >   q   �        $     Z   a         
            M     [   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  N         %   -   \      "   -   f   �   -  ��>�IJ���'�]           L      N        �   a          
          "  N      �  N           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         
     �   #   7     >   %   *   
               
        �   #   7        %   *   
                           o               n  X   l����       o         !  M     @               *  M            t   >   q   �        $  缠�p���Y췽     u   a         
            M     v   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  N         %   -   \      "   -   f   �   -           L      N        �   a          
          "  N      �  N           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7  �ݶ��⳱ϣ�     >   %   *   
                       �   #   7        %   *   
                           o               n  [   l����       o           Y   K      V      U         %  O       $         !  Q     �   >   q   �      !  O   q   �            a                #  R     �   #  S              S        
           R      Q            s              S     �   N      /   #  S     R     �   >   #  R                    O        @�Ѯ3������     s   G     �              R     �   ?      #  R     �   *  Q            Q           s   I   %  Q                          R        �      !  Q   @   4   M      #  P   !  �      q   �         !  T   q   �           -   #  U     -   L      a                  -   >   q   �           P        -   /   #  U   L      a                   !  T   q   �      !  �        U   >   q   �           ;        U   /   #  U   L      a     �=�<EMȃap�                !  2   q            #  V   !  T   q   �        U   #  P     P   L      a                     V     P   >   q           n     P   4   L        $      a         
          p  U         o               n  \   l����       o         !  M   q   �         #  V   !  2   q           n   #  P     P   L      a                     V     P   >   q   �        o     P   4   L        $      a         
            M   !  2   #  ����8�gJEg  V     n   #  P           P     :              V     P     �   4   >   #  W              P     :   	           W       3                          W     �   ?   #  W     P     �   4   #  P                                   V        P   N      p  P   K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  N         %   -   \      "   -   f   �   -           L     p�SH"Ի[�+i   N        �   a          
          "  N      �  N           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                           o               n  _   l����       o           [   K      V      U         %  O       $         !  Q     �   >   q   �      !  O  9��n(7zjb��   q   �            a                #  V     �   #  S              S        
           V      Q            s              S     �   N      /   #  S     V     �   >   #  V                    O           s   G     �              V     �   ?      #  V     �   *  Q            Q           s   I   %  Q                          V        �      !  Q   @   4   M      #  P   !  �      q   �         !  T   q   �           ��r��hU)/  {   #  U     {   L      a                  {   >   q   �           P        {   /   #  U   L      a                   !  T   q   �      !  w        U   >   q   �           ;        U   /   #  U   L      a                     X   K      V      U         %  O       $         !  Q     �   >   q   �      !  O   q   �            a                #  W     �   #  S              S        
           W      Q            s           ��C��4U�ؤ�)     S     �   N      /   #  S     W     �   >   #  W                    O           s   G     �              W     �   ?      #  W     �   *  Q            Q           s   I   %  Q                          W        �      !  Q   @   4   M      #  P   !  T   q   �         q   �           U   >   q   �           P        U   /   #  U   L      a                   !  T   q   �      !  x        U   >   q   �           �     -^����T`�     U   /   #  U   L      a                   !  T   q   �      !  �        U   >   q   �           ;        U   /   #  U   L      a                   !  2   q            #  X   !  T   q   �        U   #  P     P   L      a                     X     P   >   q           n     P   4   L        $      a         
          p  U         o               n  a   l����       o         !  M   q   �         #  X   !  2   q           n   #  2j�Ԓ�`U�  P     P   L      a                     X     P   >   q   �        o     P   4   L        $      a         
            M   !  2   #  X     n   #  P           P     :              X     P     �   4   >   #  Y              P     :   	           Y       3                          Y     �   ?   #  Y     P     �   4   #  P                                   X        P   N      p  P   K        �      ,   `         K  tW��������      *   3            �   %   -   p        =   %  �          !  �     �      %  N         %   -   \      "   -   f   �   -           L      N        �   a          
          "  N      �  N           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                        �   #   7        %   *   
                     >I�� D�<g�         o               n  d   l����       o         !  M     �               *  M            F   >   q   �        $     p   a         
            M     -   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  N         %   -   \      "   -   f   �   -           L      N        �   a          
          "  N      �  N           L      N        �   a          �
�w� �3��   
          c  �                      *   
      %   *            ,   `          �            �         !     �   #   7     >   %   *   
         "      !        �   #   7        %   *   
         "                  o               n  e   l����       o         !  	   #  Z      '      !  E   #  X     Z         (        X     ;   N      K      K      *  E             %      %        X      E          K      K        Y   K      K     !�'ǅ�
,����   	      $      &      &      #      !  
   #  Z      '      )        X         E          K           /   K      K      *  E             %      &            o               n  f   l����       o           �   K        E   K      K         1     !   K               o                  *   n  g   l����       o         !  M     �               *  M            �   >   q   �        $     �   a         
            M     ;   N      K  "�V!��zK��S      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  N         %   -   \      "   -   f   �   -           L      N        �   a          
          "  N      �  N           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         +     �   #   7     >   %   *   
         ,      +        �   #   7  # C^G��Α�        %   *   
         ,                  o                  *      n  h   l����         �   #  �   n  i   l����       o         "  Z         E   K      #  #           #     �   L      N      	      -     #     �   K      	      .      -        �   L      N      #  #      .              #   M      L        �   4     �   �   N      A         Z          K      V      =              U         %  O       $         !  Q     �   >   q  $��W&U�L��   �      !  O   q   �            a                #  X     �   #  S      /        S        
      0     X      Q            s         0     S     �   N      /   #  S     X     �   >   #  X      /      0        O           s   G     �         1     X     �   ?      #  X     �   *  Q            Q           s   I   %  Q            1              X        �      !  Q   @   4   M      #  P   !  w      q   �         !  T   q  %�����li!   �           ;   #  U     ;   L      a                  ;   >   q   �           P        ;   /   #  U   L      a                   !  T   q   �      !  }        U   >   q   �           �        U   /   #  U   L      a                   !  2   q            #  Y   !  T   q   �        U   #  P     P   L      a                     Y     P   >   q           n     P   4   L        $      a         
          p  U         o        &��m�HcM�de         n  j   l����       o         !  M   q   �         #  Y   !  2   q           n   #  P     P   L      a                     Y     P   >   q   �        o     P   4   L        $      a         
            M   !  2   #  Y     n   #  P           P     :         4     Y     P     �   4   >   #  [      2        P     :   	      3     [       3                     3     [     �   ?   #  [     P     �   4   #  P      2     '��T�
�O�*�   3         4              Y        P   N      p  P   K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  N         %   -   \      "   -   f   �   -           L      N        �   a          
          "  N      �  N           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         5     �   #   7  (�� ;+�1��#     >   %   *   
         6      5        �   #   7        %   *   
         6                  o               n  k   l����          #      $      n  k   l����       n  m   l����       o         !  M     ?               *  M            O   >   q   �        $     Z   a         
            M     [   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  N        )ͨ��]3G<Xޚ   %   -   \      "   -   f   �   -           L      N        �   a          
          "  N      �  N           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         7     �   #   7     >   %   *   
         8      7        �   #   7        %   *   
         8                  o               n  n   l����       o         !  M     >               *  M      *�6H�vfҫ��2        O   >   q   �        $     Z   a         
            M     [   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  N         %   -   \      "   -   f   �   -           L      N        �   a          
          "  N      �  N           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �         +��`T�*+0�     �         9     �   #   7     >   %   *   
         :      9        �   #   7        %   *   
         :                  o               n  o   l����       o         !  M     =               *  M            F   >   q   �        $     p   a         
            M     -   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  N         %   -   \      "   -  ,�>��oQv���|   f   �   -           L      N        �   a          
          "  N      �  N           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         ;     �   #   7     >   %   *   
         <      ;        �   #   7        %   *   
         <                  o                              n  r   l����         �   #  �      =   o         o                 -A�֙��Ak��   !  K     �   >   �  K           L      N        �   a          
          !  K     �   >   �  K           L      N        �   a          
          !  K     �   >   �  K           L      N        �   a          
          !   /   %  K            �   %  K   n        �   %  L          !  L   %  K            �   %  K   P           %  K         !   /   %  N            �   #  E   !  2   q           M   L      N           a         .�)��6E�3&�X�   
                                  =         e  �   f  �   j  �   j  �   j  �     �     �                 %   .        c                                            ]     �                             �   #  ]            n  w   l����         �   #  �   o         o         o         o         o         n  �   l����       o           �   L      N      K      K      #  �         o               n  �   l����       o        /�b�,5$���M�v   !  _     <               *  _            �   >   q   �        $     �   a         
            _     6   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  `         %   -   \      "   -   f   �   -           L      N        �   a          
          "  `      �  `           L      N        �   a          
          c  �                      *   
      %  0^S�1U�pD3zRW   *            ,   `          �            �              �   #   7     >   %   *   
         	              �   #   7        %   *   
         	                  o               n  �   l����       o           �   K      K        "   K      /   V      U         %  a       %         !  c     �   >   q   �      !  a   q   �        �   a                #  d     �   #  e      
        e     �   
           d      c            s     1�!w�x���           e     �   N      /   #  e     d     �   >   #  d      
              a           s   G     �              d     �   ?      #  d     �   *  c            c           s   I   %  c                          d        �      !  c   @   4   M      #  b   !  �      q   �         !  f   q   �           �   #  g     �   L      a                  �   >   q   �           b        �   /   #  g   L      a                  2s�浤����   !  f   q   �      !  �        g   >   q   �           ;        g   /   #  g   L      a                   !  3   q            #  h   !  f   q   �        g   #  b     b   L      a                     h     b   >   q           n     b   4   L        $      a         
          p  g         o               n  �   l����       o         !  _   q   �         #  h   !  3   q           n   #  b     b   L      a                     h  3���cg��     b   >   q   �        o     b   4   L        $      a         
            _   !  3   #  h     n   #  b           b     :              h     b     �   4   >   #  i              b     :   	           i       3                          i     �   ?   #  i     b     �   4   #  b                                   h        b   N      p  b   K        �      ,   `         K      *   3            �   %   -   p        =  4�	�H�T}ދ<<�   %  �          !  �     �      %  `         %   -   \      "   -   f   �   -           L      N        �   a          
          "  `      �  `           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                           o               n  �   l����       o  5�ڄ��/f��D         !  3     ;               *  3       &     �   >   q           $     �   a         
                o               n  �   l����       o         !  _   q   �         #  h   !  3   q           n   #  b     b   L      a                     h     b   >   q   �        o     b   4   L        $      a         
            _   !  3   #  h     n   #  b           b     :              h     b     �   4   >   #  i           6J��4)V#W�0     b     :   	           i       3                          i     �   ?   #  i     b     �   4   #  b                                   h        b   N      p  b   K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  `         %   -   \      "   -   f   �   -           L      N        �   a          
          "  `      �  `           L      N        �   a         7���S�|�}���   
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                           o               n  �   l����       o         !     #  j            !  F   #  h     j                 h     ;   N      K      K      *  F                           h      F          K      K        �   K      K     8��t��꒡�͒   	                              !     #  j                    h         F          K           /   K      K      *  F                               o               n  �   l����       o         "  M         F   K      #  #           #     �   L      N      	           #     �   K      	                    �   L      N      #  #                    #   M      L        �   4     �   �   N      A         M          K     9��l���ņ��K�   V      =   
           U   
      %  k       '   !  k   q   �           c  l              !  k   #  h     2   #  b                     b     :   	      !     h       3                     !     h     �   >   #  h     b     �   4   #  b             !        b     :         $     h     b     �   4   >   #  i      "        b     :   	      #     i       3                     #     i     �   ?   #  i     b     �   4   #  b     :�K&�����\�2   "      #         $              h   q   �      !  ~      !  f   q   �           b   #  g     b   L      a                  b   >   q   �           3        b   /   #  g   L      a                   p  k   p  b   !  f   q   �      !  �        g   >   q   �           ;        g   /   #  g   L      a                   !  3   q            #  h   !  f   q   �        g   #  b     b   L      a                     h     b   >   q     ;��jWX���5        n     b   4   L        $      a         
          p  g         o               n  �   l����       o         !  _   q   �         #  h   !  3   q           n   #  b     b   L      a                     h     b   >   q   �        o     b   4   L        $      a         
            _   !  3   #  h     n   #  b           b     :         '     h     b     �   4   >   #  i      %        b     :   	      &     i       3  <�$&��k�D
j�                     &     i     �   ?   #  i     b     �   4   #  b      %      &         '              h        b   N      p  b   K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  `         %   -   \      "   -   f   �   -           L      N        �   a          
          "  `      �  `           L      N        �   a          
          c  �                     =�"a:א�ɚ7��   *   
      %   *            ,   `          �            �         (     �   #   7     >   %   *   
         )      (        �   #   7        %   *   
         )                  o               n  �   l����                      n  �   l����                      n  �   l����         �   #  �      *   o         o                  !  ^     �   >   �  ^           L      N        �   a          
          !  ^     �   >   �  ^        >Q�e{��Gs�~     L      N        �   a          
          !  ^     �   >   �  ^           L      N        �   a          
          !   /   %  ^            �   %  ^   n           %  ^   P           %  ^         !   /   %  `            �   #  F   !  3   q           M   L      N           a          
                                  *         e  �   f  �   j  �   j  �   j  �     �     �                 %   .        c                    ?ح�Q���vm�n+                          n     �                             �   #  n            n  �   l����         �   #  �   o         o         o         o         o         n  �   l����       o         !  q     :               *  q            W   >   q   �        $     X   a         
            q     Y   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  r  @ q��`�E%0         %   -   \      "   -   f   �   -           L      N        �   a          
          "  r      �  r           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
         	              �   #   7        %   *   
         	                  o               n  �   l����       o         !  q     9               *  A�`��fn�����  q            O   >   q   �        $     Z   a         
            q     [   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  r         %   -   \      "   -   f   �   -           L      N        �   a          
          "  r      �  r           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �  B"��h�Tg�P�f�            �         
     �   #   7     >   %   *   
               
        �   #   7        %   *   
                           o               n  �   l����       o           �   K      K        "   K      /   V      U         %  s       %         !  u     �   >   q   �      !  s   q   �        �   a                #  v     �   #  w              w     �   
           v      u            s              w     �   N      /  C{'��*��մ~Q�   #  w     v     �   >   #  v                    s           s   G     �              v     �   ?      #  v     �   *  u            u           s   I   %  u                          v        �      !  u   @   4   M      #  t   !  �      q   �         !  x   q   �           V   #  y     V   L      a                  V   >   q   �           t        V   /   #  y   L      a                   !  x   q   �      !  �        D���w{�8 n  y   >   q   �           ;        y   /   #  y   L      a                   !  4   q             #  z   !  x   q   �        y   #  t     t   L      a                     z     t   >   q            n     t   4   L        $      a         
          p  y         o               n  �   l����       o         !  q   q   �         #  z   !  4   q            n   #  t     t   L      a                     z     t   >   q   �        o     E���e�	$�'  t   4   L        $      a         
            q   !  4   #  z     n   #  t           t     :              z     t     �   4   >   #  {              t     :   	           {       3                          {     �   ?   #  {     t     �   4   #  t                                   z        t   N      p  t   K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �     F��0?Y�>k�W3   %  r         %   -   \      "   -   f   �   -           L      N        �   a          
          "  r      �  r           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                           o               n  �   l����       o         !  q     8           G�Es��9�\y      *  q            w   >   q   �        $     x   a         
            q     )   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  r         %   -   \      "   -   f   �   -           L      N        �   a          
          "  r      �  r           L      N        �   a          
          c  �                      *   
      %   *            ,   `     HӍ���Lϭ       �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                           o               n  �   l����       o         !  q     7               *  q            w   >   q   �        $     x   a         
            q     )   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  r         %   -  IU�[��Rq��    \      "   -   f   �   -           L      N        �   a          
          "  r      �  r           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                           o               n  �   l����       o         !  q     6               *  q            J��8=�]?����  O   >   q   �        $     Z   a         
            q     [   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  r         %   -   \      "   -   f   �   -           L      N        �   a          
          "  r      �  r           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �  K���Ċ�b�              �   #   7     >   %   *   
                       �   #   7        %   *   
                           o               n  �   l����       o         !  q     5               *  q               >   q   �        $     |   a         
            q     2   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  r         %   -   \      "   -   f   �  L9�at�t!��q   -           L      N        �   a          
          "  r      �  r           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                           o               n  �   l����       o           �   V   
   U   
      %  |       '         !  }     �   >   q  M��ۇy�����-   �      !  |   q   �        H   a                #  z     �   #  w              w     R   
           z      }            s              w     �   N      /   #  w     z     �   >   #  z                    |   	        s   G     �              z     �   ?      #  z     �   *  }            }   
        s   I   %  }   
                       z        �      !  }   @   4   M      #  t   q   �      !  �      !  x   q   �  N�7��i��^	��           t   #  y     t   L      a                  t   >   q   �           ;        t   /   #  y   L      a                   p  }   p  t   !  4   q             #  {   !  x   q   �        y   #  t     t   L      a                     {     t   >   q            n     t   4   L        $      a         
          p  y         o               n  �   l����       o         !  q   q   �         #  {   !  4   q            n   #  t     O�V3J
��;"��  t   L      a                     {     t   >   q   �        o     t   4   L        $      a         
            q   !  4   #  {     n   #  t           t     :         !     {     t     �   4   >   #  ~              t     :   	            ~       3                           ~     �   ?   #  ~     t     �   4   #  t                      !              {        t   N      p  t   K        �      ,   `         K      *  P*�٢�J�K�   3            �   %   -   p        =   %  �          !  �     �      %  r         %   -   \      "   -   f   �   -           L      N        �   a          
          "  r      �  r           L      N        �   a          
          c  �                      *   
      %   *            ,   `          �            �         "     �   #   7     >   %   *   
         #      "        �   #   7        %   *   
         #                 Q~ߤ�wQW`���   o               n  �   l����       o         !  q     4               *  q            T   >   q   �        $     U   a         
            q     6   N      K      K        �      ,   `         K      *   3            �   %   -   p        =   %  �          !  �     �      %  r         %   -   \      "   -   f   �   -           L      N        �   a          
          "  r      �  r           L      N        �   a          
      R�Q��f�c�^      c  �                      *   
      %   *            ,   `          �            �         $     �   #   7     >   %   *   
         %      $        �   #   7        %   *   
         %                  o                              n  �   l����         �   #  �      &   o         o                  !  o     �   >   �  o           L      N        �   a          
          !  o     �   >   �  o           L      N        S)\L�	�j��6�  �   a          
          !  o     �   >   �  o           L      N        �   a          
          !   /   %  o            �   %  o   n        �   %  p          !  p   %  o            w   %  o   P           %  o         !   /   %  r          !  4   q            M   L      N           a          
                                  &         e  �   f  *   j  �   j  �   j  �     �     �                 %   .        c             T�F��N��Φ	�                                 �     �                             �   #  �            n  �   l����         �   #  �   o         o         o         o         o         n  �   l����       o           ?   K      K      K        �      ,   `         K      *   3            �   %   -   p        �   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �  U�OU+"b�s��;<      �  �           L      N        �   a          
          c  )             K               *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
         	              �   #   7        %   *   
         	              ?   K               o                  
   n  �   l����       o           �      ,   `         K      *   3            �   %   -   p        �   %  �          !  �     VN�B������Ai  �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  C                 �          #  �            *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                     !  �   !  �   q   �         !  �   q   �        W&��3��r&��H     @   a                  A   >   q   �           B   a                   !  �   q             3          #  9   p  �         o               n  �   l����       o         !  �     �               *  �            F   >   q   �        $     G   a         
          !  �   !  �     �               *  �               >   q   �        $     H   a         
          !  �   !  �     w               *  �            �   >   q   �     X۲^/��E��+     $     I   a         
          !  �   !  9   q   #        �      ,   `         K      *   3            �   %   -   p           %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  w                      *   
      %   *            ,   `          �            �              �   #   7     Y=+���2t���
  >   %   *   
                       �   #   7        %   *   
                     p  �   p  �   p  �         o                  
      n  �   l����         �   #  �                  n  �   l����         �   #  �         o         o                  !  �     �   >   �  �           L      N        �   a          
          !  �     �   >   �  �           L      N        �   a          
          !  �     �   >   �  �        Z���jRT��O�ٝ     L      N        �   a          
          !   /   %  �            �   %  �   n        �   %  �          !  �   %  �            w   %  �   P           %  �         !   /   %  �          !  9   q   #        M   L      N           a          
                                           e  *   f  H   j  �   j  �   j  �     �     �                 %   .        c                                            �     �           [?D�o8�~u��                    �   #  �            n  �   l����         �   #  �   o         o         o         o         o         n  �   l����       o         !  I   q   .        �   V   
   =   	           W      K      %  �          !  �   q   �      !  �     �               *  �            W   >   q   �        $     %   a         
          !  �   !  �     �               *  �            �   >   q   �        $     �   a         
         \�"o�_ypn9r�   !  �   !  �     w               *  �            �   >   q   �        $     K   a         
          !  �   !  p   q   @        �      ,   `         K      *   3            �   %   -   p              �          %   -   \        �          %   -   f         -   \      %  �            -   f      %  �           �                   �   %  �      (   !  �   !  �   a  �                             �            #     !     q   @  ]�Um��R��
�               #     !              #     !              #     !              #     !     q   �               #     !     q   .                        b  q               *   
      %   *            ,   `          �            �         	     �   #   7     >   %   *   
         
      	        �   #   7        %   *   
         
            p  �   p  �   p  �   p  �         o               n  �   l����       o         !  ^M��Yy ����     #  �            "  �       #  �     �                 �     :   L      L      *  �       )                    �      �       )   L      L        �   L      	                              !     #  �                    �         �       )   L        �   /   L      L      *  �       )                        o               n  �   l����       o           �       )   L      L        ;   L      /   N      #  �   !       �  _�
�?�'�� < �      #  �           �     �   N                 �     "   
                    �   !  �      c                                    4     "   K                  /   #  �           �     �   N                 �     !   
                    �   !  �      c                               M      #  �   >   q   I         #  �   !  �   q   O              �     ;              �   #  �                    ;   #  �     `�2����7�Nx�                 �   #  �     �   L      a                     �     �   >   q   I        �     �   4   L        $      a         
          p  �         o               n  �   l����                      n  �   l����       n  �   l����       o           I  t      V   	   =   
           W      K      %  �          !  �   q   �        :   N      K      K      %  �          !  �   q   �      !     q   I        �   N      K      K      %  a�S5O]�@Wg�  �          !  �   q   �        J   N      K      K      %  �          !  �   q   �        :   N      K      K      %  �          !  �   q   �        :   N      K      K      %  �          !  �   q   �        �   N      K      K      %  �          !  �   q   �      !  ~   q   H      !  N   q   2      !  O   q   3      !  =   q   &        �      ,   `         K      *   3            �   %   -   p              �          %   -   \        �      b�)�1pj�'rf��      %   -   f         -   \      %  �            -   f      %  �           �                   �   %  �      (   !  �   !  �   a  �                             �            #     !     q   &               #     !     q   3               #     !     q   2               #     !     q   H               #     !     q   �               #     !     q   �               #     !     q   �               #     !     q  c�n�;-�Vy@�Z   �               #     !     q   �               #     !     q   I               #     !     q   �               #     !     q   �                        b  (               *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                     p  �   p  �   p  �   p  �   p  �   p  �   p  �         o               n  �   l  d��6C��3������       o           ~   h     �   #  �         o                                    n  �   l����         �   #  �     �     �              �   !  �      c                               o         o                       #  �   !  �     �   >   �  �           L      N        �   a          
          !  �     �   >   �  �           L      N        �   a          
          !  �     �   >   �  �           L      N     e�yC³��`P�     �   a          
          !   /   %  �            �   %  �   n        �   %  �          !  �   %  �            #   %  �   P           %  �         !   /   %  �          !  I   q   .        M   L      N           a          
          !  ~   q   H        �   L      N           a          
          !     q   I        �   L      N           a          
               #  N        #  O   !  =   q   &        M   L      N          fhp�k�';Ak   a          
            �   #  �                                    e  H   f  C   j  �   j  �   j  �     �     �                 %   .        c                                            �     �                             �   #  �            n     l����         �   #  �   o         o         o         o         o         n     l����       o           �      ,   `         K      *   3            �   %   -   p        g:����<�{�M  �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  D                        *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
         	              �   #   7        %   *   
         	            #  <         o               n  	   l����       o           <      h�s�x��)��R  ;          V   
   =   
           #  �   !  �   q   �        H   !  �   q   �        H   !  �     K   a  �      �       !  �   #  �     2   #  �            
        �     :   	           �       3                          �     �   >   #  �     �     �   4   #  �      
              �     :              �     �     �   4   >   #  �              �     :   	           �       3                          �     �   ?   #  iM��"�w��  �     �     �   4   #  �                                   �   q   �      !  v      !  �   q   �           �   #  �     �   L      a                  �   >   q   �           [        �   /   #  �   L      a                   p  �   p  �     <      ;          K      K      K        �      ,   `         K      *   3            �   %   -   p        �   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -     j��w2�0g!8$T:        L      N        �   a          
          "  �      �  �           L      N        �   a          
          c  {                      *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                       :   #  �   #  �                    �     �   
           �     �   >       3                          �     �  ky�¿���	;�Y   /   #  �                          �   q         !  �   q   �              �   >   q   �           �     �   4     �   #  �   #  �           �     �              �   #  �                    �        �   /   #  �   L      a                   !  �   q   �         #  �   !  �   q   �              n     �              n   #  �                    �   #  �                    �   #  �     �   L      a                  lZ��{�q9���,     �     �   >   q   �        n     �   4   L        $      a         
            �   h     �   #  �   p  �         o                                    n     l����         �   #  �     �     �              �   !  �      c                               o         o                       #  �   !  �     �   >   �  �           L      N        �   a          
          !  �     �   >   �  �           L      N        mg�5�&)��^hƝ  �   a          
          !  �     �   >   �  �           L      N        �   a          
          !   /   %  �            �   %  �   n           %  �   P           %  �         !   /   %  �            �   #  <                                    e  C   f  w   j  �   j  �   j  �   g     g      g   �   g   �     �     �                 %   .        c                                            �     �                    n�;�,�0��9D�           �   #  �            n     l����         �   #  �   o         o         o         o         o         n  (   l����       o         !  w      �   q                  #  �        E   a                #  �           �     �         	     "   #  �            	        �   q             3         !         3                
     "   #  �            
        !   #  �                             �         o           ox2BR	�;�x�            n  )   l����       o         !  G   q   -         #  �      �   q           -   #  �     �   L      a                         o               n  *   l����       o         !  :   q   $         #  �      �   q           n   #  �     �   L      a                         o               n  +   l����                      n  +   l����         �   #  �   n  ,   l����       o         !  �        q                  #  �        p��E��\S��x  7   a                #  �           �     �              !   #  �                    �   q             3         !         3                     "   #  �                    !   #  �                             �         o                     n  -   l����       o           �   #  G         o               n  .   l����       o               #  �     4   #  �           �     :              �     �     �   4   >  q�j34+r<@Bt�   #  �              �     :   	           �       3                          �     �   ?   #  �     �     �   4   #  �                                   �   !  �      q            !  �   q   �           V   #  �     V   L      a                  V   >   q   �           �        V   /   #  �   L      a                   !  �   q   �      !  v        �   >   q   �           [        �   /   #  �   L      a               r��*�O����(      !  �   q   �         �   q              �   >   q   �           n        �   /   #  �   L      a                   !  :   q   $         #  �   !  �   q   �              n     �              n   #  �                    �   #  �                    �   #  �     �   L      a                     �     �   >   q   $        n     �   4   L        $      a         
          p  �         o               n  /   l����         s���T��*�Y               n  /   l����         �   #  �   n  0   l����       o         !  :   q   $         #  �      �   q           n   #  �     �   L      a                         o                        n  1   l����         �   #  �            n  2   l����         �   #  �   n  4   l����       o         !  G   q   -      !  �     �               *  �            �   >   q   �        $     I   a         
          !  �   !  :   q   $        t0�kxoJ|Ň
�  �   V   
   =   	           W      K      %  �          !  �   q   �           q         !  �     �               *  �            F   >   q   �        $     �   a         
          !  �     ;   X      =   	           W      K      %  �          !  �   q   �      !  �     w               *  �            �   >   q   �        $     G   a         
          !  �   !  p   q   @        �      ,   `         K      *   3            �   %   -  u��>�|�7�WdQ@   p              �          %   -   \        �          %   -   f         -   \      %  �            -   f      %  �           �                   �   %  �      (   !  �   !  �   a  �                             �      
      #     !     q   @         	      #     !        	      #     !     q   �         	      #     !        	      #      !      q            	      #  !   !  !   q   �         	      #  "   !  "   q   $  v�6�-�"�装2          	      #  #   !  #      	      #  $   !  $   q   -         	         
   	   b  n   	            *   
      %   *            ,   `          �            �              �   #   7     >   %   *   
                       �   #   7        %   *   
                     p  �   p  �   p  �   p  �   p  �         o                              n  8   l����         �   #  �         o         o                  !  �     �   >   �  wm{1P?�옹H  �           L      N        �   a          
          !  �     �   >   �  �           L      N        �   a          
          !  �     �   >   �  �           L      N        �   a          
          !   /   %  �            �   %  �   n           %  �   P           %  �         !   /   %  �          !  G   q   -        M   L      N        %   a          
          !  :   q   $        M   L      N           a          
         x�|�Q6����u�{                                    e  w   f      j  �   j  �   j  �   g     g     g     g     g     g     g     g     g     g     g     g  	   g     g     g     o         o         o         o         j  �   l����          .        #  �     �   %   .          �   %   -   Y        �     �              �     =              �             9     �   %   -   Y         \     9        �     �        :     �   %  y�y���5ᰐ�   -   Y         �      s  E  E   !   H   !  &   *   H       "     6   s  �  �   !  �   !  &   *  �       "     7   s  %  %   !   H   !  &   *   H       "      �           ;        �   %   -   Y        8     :        �     �                        -   H        �        <      ,   `        �   *   3          !   /     �   c  �                <        �   %   W   �   !   !  '   #  �     4     =           #           #          #  zZ..wB"�&���]          #          #          #          #          #          #          #          #       	   #  
        #          #          #        -   [        �        >     �   %   /   �         \      !  (   #  �     3     ?      !   /   c  �                >         -   Y        �        @   j  �   l����       m       �   a  �       �           3              3             V      U         %   *   $   *   #  6  {�1�\m	He�oM     A   k  �   l����         B        �   #  6     �   %   *   $   *     A        6   V      U         %   *   $   *     @      k  �   l����       j  �   j  �   j  �   l����       n BA   o           �   %   -   H         -   [        �        C   !  �   %   /   �      !  �      %  �   0      %  �   @        �      %  �   	      %  �  �      !  )   %  �   �   "     C        �   #  �      -   Y        �        D     �   %   -   Y        |� �=N{�����  �   %   -   H        8     D      !   *     *   >   q   =           L      N        +   a          
          !   *     ,   >   q   =           L      N        �   a          
          !   *     -   >   q   =        s   L      N           a          
             -   [        �        E     �   %   -   [         	     F     E        �     �         
     F         	           %   *            
        	   %   *           �  }
�+"*`�V�   #   6     �   %   W      !      W   m   !     �         i   "   W   d   q   P        �   L      N        .   a          
                   i      "   W   d   q   P        �   L      N        .   a          
             W   �   !     �         j        %   /   �               j        �   %   W   �   !           �               W   m   !     �              �   #               X         /   �        �   
     G      /   �        �  ~ZwS����+�
�        H      /   �          2   �   "             I      /   �          2   �      !  /   *   2       "      /   �          2   �   "        I         5        H        G         /   �      #   7   j  �   l����          /   �          2   �   "   %   .   p   "      /   �          2   �   "             J      /   �          2   �      !  0   *   2       "     J      c                  k  �   l����          5         Y         /   �      #   7   !   /  ��]#��8�ʹ        c  �                                  %   *                     W   m   !     �                 %   *                 6      n   �   l����         �  �        �        L   !  �       3          %  �   %      "   W       %  �   �      !  1   %  �   `   "     �   %  �  �        K     5        �   0          3          #  �   n   �   l����       !  >     �     �   >       3          *  >          n   �   l����       !  L     �  �P�d�PPG���     �   >       3       +   *  L       +      H        L        �   %  �   
        �      #   7   %   /   �         /   �        �   	     M     �          %   *   �        �  �      %   *   �        �   
       %   *   �         �   L      %   *  c        M         /   �      #   7   j  �   l����            %   .   p   "   c                  k  �   l����         K         H                    %   *         n   �   l����       o           �  �(�_��7�W}�      ,   `         K      *   3            �   %   -   p        �   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
                j  �   l����       j  �   j  �   l����             c  v                   k  �   l����       k  �   k  �   l����          *   
      %   *            ,   `          �            �dA��ɩ:n�|  �        N     �   #   7     >   %   *   
        O     N        �   #   7        %   *   
        O                  o               n   �   l����       o                 j       ,     �      ,   `         K      *   3            �   %   -   p        �   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a  ��	�t,���ї�}          
                j  �   l����       j  �   j  �   l����             c  -                   k  �   l����       k  �   k  �   l����          *   
      %   *            ,   `          �            �        P     �   #   7     >   %   *   
        Q     P        �   #   7        %   *   
        Q                  o               n   �   l����       o           �      ,   `         K      *   3            �   %   -   p        �   %  ���F���L��  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
                j  �   l����       j  �   j  �   l����             c  H                 �       -   #  �         k  �   l����       k  �   k  �   l����          *   
      %   *            ,   `          �            �        R     �   #   7     >   %   *   
     �k���Xj�w�E�     S     R        �   #   7        %   *   
        S            !  }   q   G         #  �   !  �   q   �        �   #  �     �   L      a                   p  �         o               n   �   l����       o         !  �            _                      *  �               >   q   �        $     �   a         
            �     �      ,   `         K      *   3            �   %   -   p        �   %  �          !  �     �     �4� m,��&`~�   %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
                j  �   l����       j  �   j  �   l����             c  �                   k  �   l����       k  �   k  �   l����          *   
      %   *            ,   `          �            �        T     �   #   7     >   %   *   
        U     T        �   #   7        %   *   
  ����ooyn��N        U                  o               n   �   l����       o           �      ,   `         K      *   3            �   %   -   p        �   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
                j  �   l����       j  �   j  �   l����             c  �                   k  �   l����       k  ��+xsU����6�  �   k  �   l����          *   
      %   *            ,   `          �            �        V     �   #   7     >   %   *   
        W     V        �   #   7        %   *   
        W                  o               n   �   l����       o           �      ,   `         K      *   3            �   %   -   p        �   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
  �Ͽ��R.����          "  �      �  �           L      N        �   a          
                j  �   l����       j  �   j  �   l����             c  �                   k  �   l����       k  �   k  �   l����          *   
      %   *            ,   `          �            �        X     �   #   7     >   %   *   
        Y     X        �   #   7        %   *   
        Y                  o               n   �   l����       o           �      ,   `  �v+d#���ړ���         K      *   3            �   %   -   p        �   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
                j  �   l����       j  �   j  �   l����             c  �                   k  �   l����       k  �   k  �   l����          *   
      %   *            ,   `          �            �        �����L; ̸  Z     �   #   7     >   %   *   
        [     Z        �   #   7        %   *   
        [                  o               n   �   l����       o           �      ,   `         K      *   3            �   %   -   p        �   %  �          !  �     �      %  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
                j  �  ��������0   l����       j  �   j  �   l����             c  �                   k  �   l����       k  �   k  �   l����          *   
      %   *            ,   `          �            �        \     �   #   7     >   %   *   
        ]     \        �   #   7        %   *   
        ]                  o               n   �   l����       o           �      ,   `         K      *   3            �   %   -   p        �   %  �          !  �     �      %  ��e�'��Ri�S  �         %   -   \      "   -   f   �   -           L      N        �   a          
          "  �      �  �           L      N        �   a          
                j  �   l����       j  �   j  �   l����             c  *                   k  �   l����       k  �   k  �   l����          *   
      %   *            ,   `          �            �        ^     �   #   7     >   %   *   
        _     ^        �   #   7        %   *   
     �qŰHf��'�Q�     _                  o               n   �   l����       o              #   �         o               n   �   l����       o               o                     l����          	              
   %   *         l����               7        �  �        �        c     �   %  �   
        #      #   7   %   /   �         /   �        �   	     d     �          %   *   �        �  �      %   *   �        �   
       %   *   �         �m����	f�$��  �   L      %   *  c        d        `     c        �  �        �   �           b     �   0          3   0      %  �  �        �         %  �   0        b        �             3           �   	     a     �                      3                 3         K      >   *   3                 3         K           4   K      *   3           �   %  �  �        `     `     a      j  �   l����       !   /   !   R   q         c  �  ��J���*�r*�E              k  �   l����         `        �         Z      c                     5               j  �   l����          W   m   !     �        e           f     e              f                 =   %   /   �                     !  2   #  �     1     g      !  3   #  �     .     h                  /   �        �   	     i     O      /   �           j     �      7        j   !   /     �   c  �                k     j     �n���:�P�h�   !   /     �   c  �                k        l     i        �   %   -   H         W   m   !     �        m     �   %   /   �        �   %   -   [        n     m        �   %   /   �        �   %   -   [        n         /   �         ,   `         K      *   3            l            k  �   l����       j  �   l����         1        �      k  �   l����       j  �   l����         3        s   %  #          !  �   %  �               %  ���d:L~�-���  �         !  �   %  �               %  �   0           %  �   @           %  �   P           %  �   `   "        %  �   p   "        %  �   �           %  �   �   "        %  �   �   "        %  �   �   "        %  �   �           %  �   �           %  �   �           %  �              %  �             %  �  0           %  �  p   .        %  �         !  �   %  �               #   !        %   *       /   !  ����NL;#��   *     4   >   q   =        M   L      N        5   a          
               #           #           #        s   #         s   #   "        #   7        %   -   q           %   -   r      !   -     6   >   �   -        M   L      N        �   a          
          !   -     7   >   �   -        M   L      N        �   a          
          !  8   %   .       "   !  9   %   .   �   "   !  :   %   .   �   "        %   /   �           %  �1#�>���x��   /   �           %   /   �      !   W   q   P        s   L      N        ;   a          
               %   W           �   %  �       0     �   #   (     �   #  +     M   #  >        #  ?   !  A   q   *        M   L      N        -   a          
            �   #  J   !  L   q   0        M   L      N        <   a          
            �   #  M     �   #  S     W   #  T     $   #  U     =   #  V     �   #  X     �   #  Y     �  �|{<�k�<d�[ܗ   #  Z     �   #  [     �   #  b   !  o   q   ?        M   L      N        6   a          
          !  p   q   @        M   L      N        �   a          
               #  t     �   #  u   !  }   q   G        M   L      N           a          
            �   #  �     �   #        �   #  �     �   #  �     �   #  �        #  �        #  �        #  �        #  �        #  �     �      k  �   l����       j  �   l����      ���z���1�JI7     4        �      k  �   l����       j  �   l����         .        �   %  �   
         �  �        �        o   !  �   %   /   �        �   %   /   �      j     l����       !   /     �        #  #   c                k     l����       !  �      %  �   0      %  �   @         /   �        �   
     p      /   �      #   7   j  �   l����            %   .   p   "   c                  k  �   l����         p        o        �      k  �   l  ���z=#찻����       k  �   l����       k  �   k  �   o         o         j  �   l����         /        �   %  �   
         �  �        �        q   !  �   %   /   �        �   %   /   �      j     l����       !   /     �        #  #   c                k     l����       !  �      %  �   0      %  �   @        q        �      k  �   l����                j  �   l����         �   %   -   [      !  =   #  �     /     r         /   �        O        ��CA���q�@+  s      ,   `        �   *   3            t     s         ,   `        �   *   3            t         [   k  �   l����                n BB      7   #   7      [        8        u     u         e      f  �   j  �   j  �   j  �   g  �      .          T              �   %   .                       c                    �   %   -   H        �   %   -   [                        e  �   f      j  �   j  �   j  �   !   /      7   c  �  �r
�����\J                                e      f      j  �   j  �   j  >   j  A     �   #  ?     �   a          �       %  ?           C     B   a          �         �   a                 a          �             c  D                        a  �              #  �     �   #  �              �     K              �     �   
         !  �     �   A           *  �                         !  �     �   A        �     �   /   a  �            ��}$�eڅݐ��       3          *  �                     �     �   /   #  �                    �            �           �            �   0        �   @        �   P        �   `        �   p        �   �        �   �        �   �        �   �        �   �        �   �        �   �        �   #  �     �   %  �       1   !  �   c                                 F   a           �       !  ?   c  G                 e             l      q      �8_�\�5���v  �          `     �      �   `           �      �   p      `     V      �   �      
     �      �   �           �      �               �      �  @           �      �  P           �      �  `           �      �             �       +   P           �      �               �      �               �       +   0            W       +   @            7       +   �           �       +   �           �       +   `           �       +   �  �ه�-�"E���/           �       +               �       +   �           �       +   �           �       +   �           �       +   �           �       +   �      
     �       +   �           �       +   �           �       +   �           �       +   �           �       ,   �           �       ,   �           �       ,   �           �       ,   0           �       ,   �           �       ,  
           �       ,   �           �       ,   �        ��9ˏ�&����m     �       ,   �           �       ,   �         
  �       -   H           �       -   [           �       -   Z           �       -   V           �       -   0           �       -   L         
  �       .                     .                     .                    .                    /   0            +       /   @            ,       /   P            -       /   `            .       /   �            0       /   p            *  �E�D�9��U���@       /   �                  /   �                  /   �         
  	      �          �     
      �          �     �      �                	
      �          
     	*      �               	4      �               	5      �               	6      �               	7                     	8                      	9      9               	:      J               	;      ]               	<      n               	=      �               	>      �  ����ʑ5�ͺ�ߔ               	?      �               	@      �               	A       ,  	           	B       /               	B      �                /       '               	C      �               	G      �               	e      �               	�      �               	�      �               	�      �               	�      �               	�      �               
      �          
     
7      �          
     
A      �          
     
K      �         �׬�^c��]�"   
     
U      �          
     
_      �          
     
i      �          
     
s      �          
     
}      �          
     
�      �          
     
�      �          
     
�      �          
     
�      �          
     
�      �          
     
�      �          
     
�      �          
     
�      �          
     
�      �          
     
�      �          
     
�      �          
     
�      �          
     
�      �   �            ����G�����       �   �            � <�   �   �           :�   �  �   �          ��          $                 )   "     *   +             -   ;             5   I             C   T             D   b     H   m             W   |     v   �             w   �             x   �             {   �     �   �     �   �     �   �             �   �             �               �               �  ,             �  <             �  h     �  z       �       �  �t�O��/���       �       �       �       �       �     l                                   �       �  ,     �  A     �  O             �  _     �  s     �  �     �  �     �  �     �  �     �  �     �  �     �  �     �       �          +                =      �     �  S     @  g     D  w     G  �                      ��������@@@@@@@@@@@@@@@@@@@@@@�                                                                       �Y<y��,c��hTj                                                       |   ��                                                                       ��0                                                                                                                                                                                                                                                                      �   "                                      �                              �              ��r����(�0~�   &               (                                       	      )         
      ,                              #                              +                                                                           
                                             	                                                            (                                                                    ��������"A��                         
         !      :         "                 $           @    �� ��                                                                                                                                                                                                                                                                                                                                                                                                                      ��t�V�*��c@�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   �    � [�D         ��%  !N7�        �:�3
                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ��Z4�=�8�b�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��s�Xo   �@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   �`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   �  �����                                  0                                     P  `  P ���������� @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                ��������@@�����@@@@@������@@@@@@@@@@@@@@@            \���@@@@@@@@@@@@@@@@\������@@@@@      �          @@@@@@@@@@@@@@@@@@@@@�@@@@@@@@���������������������������������������������������@@@@��������@@�������@@@@@@@@@@@@@@@@@@                                @@                     0      0          ��������@@����@@@@@@          ��5���[M��m	H  ��d�ya[OI��������@@@@����@@@@@@          ������@@@@@@@@@@������@@@@����@@@@@@          ������@@@@@@@@@@��������@@����@@@@@@          ��������@@@@@@@@������@@@@����@@@@@@           D�����9{���.���������@@����@@@@@@   :       ��������@@@@@@@@                                                                                                                                                                                                                                                                                  ���L�3����c��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��s�Xo   �`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   �   P� [�D         :�3
  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           ��:ª��*� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��s�Xo   �@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   �`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   �                                  ���@⨔���@あ��      V  �@   @  
@  p  �  
�  �            ���� � ��� ���� �� \���m�� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \����  �% ��S���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� \  ���,`S!����� \���� \���� \���� \���� \���� \���� \���� \���� \���� \���� ����� ������� ������� ����� �������� �������� ������ ��������� ��������� ������� ���������� ���������� �������� �������� ������� ������ ������ �������� ����� ������ ������ ��������@@                     ��������� ���������� ������ �������� ������ ��������� ������ ��� ������ ����������� ����� ������������ ������� ���������� ����������� � � � ������� ��������� ������� ������� ����������� ��������� m����m����m����������� �������������� � ��������  ����^+��؂;�� ������������ ������������ ����������� �������� ��������� �� �� �� ���������� ������ ������m� ��������� ������� �������� ����� ������ ����� m����m����m������� m����m����m�������� m����m����m����� m����m����m������ �������� \�� m����m����m������� m����m������m������� m����m����m���������� m����m������m���������� m����m����m����������� m����m������m����������� m����m����m����� m����m������m����� m����m����m���������� m����m������m���������� m����m����m���������� m����m������m���������� m����m����m�����������  � 1""y�ĜM1� m����m������m����������� m����m����m���������� m����m������m���������� m����m����m��������� m����m������m��������� m����m����m��������� m����m������m��������� m����m����m������ m����m������m������ m����m����m������� m����m������m������� m����m����m������� m����m������m������� m����m����m������� m����m������m������� m����m����m����� m����m������m����� ���� ���� �� ���� ���������� ���� ��������� �m�������� �m����� �m����� �m������ ���������� ������ ���������� ��������� ��������� ����� ����� ����������� �����  �x�����d�E˙�� ��������� ������� ������� ����������� ��������� ���������� ���������� ������� ���������� ���������� �m����� �m����� ��������� ��������� ������� ������� ����                           
�                       ����                  
�                      ����                                        ����                  @                       ����                  p   @                                        �                    
                        �                                   ��>Wˆ[�n��|                                  	                  0                        
                  `   0                                      �   @                                      �                                            �   �  �                                                                                P                                           �                                            �   @                	                        �                     ǈrQ�%��Q��	                                           	                        @                    	                        p   @                                        �                                            �   @                
   ����                                                              0   �   �      �                            `       	                 +                  �                       .                  �                       0                  �     ȑr��e݁~����                                                   �                            P  (  (      �                            �            �                            �              �                            �   p   p      �                                        �          "                  @   `   `      �          $                  p   P   P      �          %                  �   �   �      �          &                  �   8   8      �          '          ɍ�3���a-�             0  0      �          *                  0   �   �      �          ,                  `   0   0      �          /                  �   h   h      �          1                  �  �  �      �                            �     �               ����                                          ����                  P      �   E           ����                  �                       ����                  �      P   G           ����                  �      �             ��\�W��t8Y��      )                    @  �             ����                  @                       ����                  p         E           ����                  �                       ����                  �      p   K           ����                         �  @              (                  0  }   �  P           ����                  `                       ����                  �      0   E           ����                  �                       ����                  �      �A;P$�^9�܎�  �   P           ����                         �  `                                P    �  �          ����           S      �  �  3�  3�  0       ����          !      �   �  Q�  Q�   �       ����          F      �  �  Rp  Rp  �       ����          �        h  T   T    0       ����          �      @  �  TP  TP   0       ����          �             T�  T�   0         �                        �  T�      �                     *�      {x      �                 *�  *�  ̈��r�!zo�>   �  }                        +@  +@   �  4      4                 ,   ,    �  �l      [                 ,�  ,�     ��      �                 -�  -�   `  �       �                 .  .   �  ��      �                 .�  .�   `  �(      �   	              /0  /0   `  �      �   
              /�  /�   0  �      �                 /�  /�   0  ��      �                 /�  /�  P  ��      $                 1@  1@   `  ��      ?                 1�  1�  �  �|      �                 ��f鈊����o�'      3�      ��                                       0  !�     	T  J                           `  �  �  �                             �  �  �  �                             �  P  �  [  
                           �        �   �       ����                         P   S   W                                   �  i                             �  �  �  1                                     �  	/                                      �  		        νD��OR�l6�}�                         `  �                               @  �  �                               p  �  �  �                                     �  �                                     �  =                                0  �  �                                     �  �                                     �  �                             �  �  �  J  	                               �  �  �                                     �ָ��&�w΂�}  �  T                                P  �                                       �  	                                     �  �                             �   �  �  �  5                           �   0  �  �                               �  �  �                             @  p  �  �                                     �  �                                     �  (                             �      �  �                     Й�ºb��B E�                  �  �                                     �  �                              `   �  �  �  *                                   �  n                              �      �  �  -                                      	B  +                           !   !�  �  $  C                           !P  !�  P  	L  ?                                   �  	G  >          %                         p  	O  A                                   �  �  H      ѿ%��{š%1,��                        "  &`  0  
)            $                 "@  %  @  	�                             "p  #�     	�  Y                           "�  #0  P  	y  T          (                 "�  #      	d  M          '                         �  	_  L                                   P  	n  S                           #`  #�  P  	�  V                                   P  	�  U                                      	�  X          +                 #�  $�  �30u�~�a��9  `  	�  
                           $   $P     	�  [          )                         �  	�  Z          *                            	�         ����                 $�  $�  �  �   *          $                         @  	�             .                         �  	�            +                 %@  %�  `  	�            $                 %p  %�  @  	�                                        	�  b                                    0  	�            +         ә�d:C��	��          &   &0  `  
            /                         `  
	            0                         �  
                             &�  (  �  �  v       ����                 &�  'P  �  F  o          .                 &�  '   �  
1                                     �              0                         �  
<                             '�  '�  P  
G  t       ����                         �  !  p                           '�      �  �         ��܀Xu��                               P  
O  u                           (@  )0  �    �                           (p  (�  �  �  x                                   �  ?  w                           (�  )      
W  �                                   �    }                                      
a  �                           )`  )�  �  �  �                           )�  )�  �  [  �                                   �  4  �                                   �/���i�=v�'��  �  �  �                           *   *P     
k  �                                   �  �  �                               *�    
s  �                                   P  
{  �                           *�  +       @                                   P    7                                   �    k                           +p  +�  P  -  &                                   �  "  %                           +�      P  )  K                   ֙�JP�!�{�П                  P    8                           ,0  ,`  P  S  .                                   �  F  ,                                   �  @  �                           ,�  -   P  S  /                           ,�         r  '                                   P  f  $                           -P  -�     t  r                                   �  x  ^                                      v  s                           -�      P  �  |      ׼o��A���>�                               P  S  0                           .@  .�  P  �  y                           .p      P  S  1                                   �  �                                     P  �                             /          �  E                                   P  S  2                           /`         �  F                                   P  S  3                                   P  S  4                                   ج��v�]��U�<  P    9                           0   0�  P    N       ����                 0P        �  I          "                           !  =                           0�  0�  �    ~                                   P    O                               1  �           ����                         @  �  �                               1p  P  /  <                                   �  6  <          &                 1�  2�  �  g  G                   ٘vxX-�ؿY\ll          2   2`  �  �   �                               20  �  �                                      �  �   �                           2�  2�  P    :                                   �  m            %                         p  Q             &                 3   3P  �  Z   �                                   P  `   �          $                         @  I              �             3�  B   �   �   �            �             3�  :�  �  �  8      ��x{��[!�U��        �             4  6   �  m               �             4@  50  �    �            �             4p  5   �  �  �            �             4�  4�  �  �  x            �                     �  �  p            �                     �  �  �            �                     �    �            �             5`  5�  �  a              �             5�  5�  �    �            �                     �    �            �                     ۝�S����mC�S�  �    �            �                     �  g              �             6P  8`  �  �  �            �             6�  7p  �  �  P            �             6�  7@  �  �  @            �             6�  7  �  y  0            �                     �  s  (            �                     �    8            �                     �  �  H            �             7�  80  �  �  p            �             7�  8   �  �  `            �     ܙ��3^_�e	�                  �  �  X            �                     �  �  h            �                     �  �  x            �             8�  9�  �  �  �            �             8�  9P  �  �  �            �             8�  9   �  �  �            �                     �  �  �            �                     �  �  �            �                     �  �  �            �             9�  :@  �  �  h            �             9�  :  �  �  �      ݦD~��(�D��        �                     �  �  �            �                     �  �  �            �             :p  :�  �  �  (            �                     �  �               �                     �  �  0            �             ;   ?P  �   [               �             ;0  <�  �  +  �            �             ;`  ;�  �  �  X            �             ;�  ;�  �  �  H            �                     �  �  @            �                     ޝ��c^<��2{�  �  �  P            �             <   <�  �    �            �                 <P  �  �  `            �                     �  U               �                     �  %  �            �             <�  >0  �  �  �            �             =  =�  �  C  �            �             =@  =p  �  7  �            �                     �  1  �            �                     �  =  �            �             =�  >   �  [              �     ߘQ9m�}t���                  �  I  �            �                     �  �  �            �             >`  >�  �    �            �             >�  >�  �    �            �                     �  �  �            �                     �  	  �            �                 ?   �                 �                     �                �             ?�  @�  �   �   @            �             ?�  @  �   m                �                 ?�  �   a         ৷�4�����        �                     �   g               �             @@  @p  �   y   0            �                     �   s   (            �                     �      8            �             @�  A�  �   �   `            �             A   A`  �   �   P            �                 A0  �   �   H            �                     �  O  �            �                     �   �   X            �             A�  A�  �   �   p            �                     ᙾ�a-n�<F  �   �   h            �                     �   �   x            �             BP  K   �  �               �             B�  EP  �                 �             B�  D   �   �   �            �             B�  Cp  �   �   �            �             C  C@  �   �   �            �                     �   �   �            �                     �   �   �            �             C�  C�  �   �   �            �                     �   �   �            �     ��A��Y�QS�0                  �   �   �            �             D0  D�  �   �   �            �             D`  D�  �   �   �            �                     �   �   �            �                     �   �   �            �             D�  E   �  	   �            �                     �     �            �                     �     �            �             E�  HP  �  u  �            �             E�  G   �  E  @            �             E�  Fp  �  -         �<eD<����:��        �             F  F@  �  !              �                     �                �                     �  '              �             F�  F�  �  9  0            �                     �  3  (            �                     �  ?  8            �             G0  G�  �  ]  `            �             G`  G�  �  Q  P            �                     �  K  H            �                     �  W  X            �             G�  H   ��0�0�|�m<  �  i  p            �                     �  c  h            �                     �  o  x            �             H�  I�  �  �  �            �             H�  I@  �  �  �            �             H�  I  �  �  �            �                     �  {  �            �                     �  �  �            �             Ip  I�  �  �  �            �                     �  �  �            �                     �  �  �            �     ��b-��J����          J   J�  �  �  �            �             J0  J`  �  �  �            �                     �  �  �            �                     �  �  �            �             J�  J�  �  �  �            �                     �  �  �            �                     �  �  �            �             KP  N   �  5  �            �             K�  L�  �    @            �             K�  L@  �  �               �             K�  L  �  �        �(F P���P�*        �                     �  �              �                     �  �              �             Lp  L�  �  �  0            �                     �  �  (            �                     �  �  8            �             M   M�  �    `            �             M0  M`  �    P            �                     �    H            �                     �    X            �             M�  M�  �  )  p            �                     �<��z���?  �  #  h            �                     �  /  x            �             NP  O�  �  e  �            �             N�  O  �  M  �            �             N�  N�  �  A  �            �                     �  ;  �            �                     �  G  �            �             O@  Op  �  Y  �            �                     �  S  �            �                     �  _  �            �             O�  P`  �  }  �            �     ���`t�"�2          P   P0  �  q  �            �                     �  k  �            �                     �  w  �            �             P�  Q   �  �               �             P�  P�  �  �  �            �                     �  �  �            �                     �  �  �            �             QP  Q�  �  �              �                     �  �              �                     �  �               '�             Q�  R  0  '          �|DP�/�;�         '�                     0  /              &  '�                 R@  �  7   @            '�                     �  =   x          &  &�             R�  S`  �  j   `             &�             R�  S   0  V                 &�                     0  `   @             &�                 S0  0  }   �          1  &�                     �  �                &�             S�  S�  0  O                &�                     �  r   �             &�             S�      �U�q)�=.��^��  0  �   �             &�                     0  �   �          ,  $�                     0  �  8             0                      0  �  �            1                     �  �           e                  Xt  q|  Wx  n�  m�  ]�  q  o�  u�  v�  zX  z�  u$      s�  V�  Zl  ZH  Z�  s,  t�  vD  Y(  [D  s�  [�  ]�      y\  w@  s  nd  z  v�  p�  {T  o�  [�  w�  sP  tp  w�  XP  W�  w  n�  X�      wd  \d  z�  tL  x�  z�  ]  ]`  \�  ]�  x�  t�  r0  uH      y�          _  o<  _|  _X  u�  ����ȹj��T�  _4  _�  y�          y�  {0  z4  vh  y�  x`  z|  x�  i�  j  w�  l�  lH  m   y  x<  l�  t�  mh  m�      {      y8  u�  	T  Vl                             �  V�              0              �  V�              `              [  V�              �              �  V�              �               S  W               �               �  WD              3�              �  Wh              3�              m  W�              3�                W�              4              �  W�              4@          �<괥�lvI0�9�      �  W�              4p              �  X              4�              �  X@              4�                Xd              5               a  X�              50                X�              5`                X�              5�                X�              5�              g  Y  V�          5�              �  Y<              6               �  Y`              6P              �  Y�              6�              y  Y�              6�              s  Y�              6�                폵x�B��ʵf�  Y�              7              �  Z              7@              �  Z8              7p              �  Z\              7�              �  Z�              7�              �  Z�  V|          8               �  Z�              80              �  Z�              8`              �  [              8�              �  [4              8�              �  [X              8�              �  [|              9               �  [�              9P              �  [�              9�              �  [�  X  �OI�5�}Ewy�          9�              �  \              9�              �  \0  W�          :              �  \T              :@              �  \x              :p              �  \�              :�               [  \�              :�              +  \�  Yp          ;               �  ]              ;0              �  ],              ;`              �  ]P              ;�              �  ]t              ;�                ]�  Y�          ;�              �  ]�              <               U  ]�              ���e�[�JN���  <P              %  ^  Y�          <�              �  ^(              <�              C  ^L              <�              7  ^p  YL          =              1  ^�  Z           =@              =  ^�              =p              [  ^�  W�          =�              I  _   X,          =�              �  _$              >                 _H              >0                _l              >`              �  _�              >�              	  _�              >�                _�              >�      ���{���K#@�H�            _�              ?                �  `               ?P               m  `D              ?�               a  `h              ?�               g  `�  W          ?�               y  `�              @               s  `�              @@                 `�  W0          @p               �  a  `x          @�               �  a@  \�          @�               �  ad              A               O  a�  ]<          A0               �  a�  `T          A`               �  a�  `�          A�              �
�V!��g�˸   �  a�  `0          A�               �  b  `�          A�              �  b<              B                 b`  a�          BP               �  b�  b          B�               �  b�  a�          B�               �  b�  aP          B�               �  b�  `          C               �  c  b(          C@               �  c8  a�          Cp               �  c\  a          C�               �  c�  bL          C�               �  c�  c           D                �  c�  b�          D0               �  c�  �K7�0mh�y��  `�          D`               �  d  b�          D�              	  d4  cH          D�                dX              D�                d|  c$          E               u  d�              EP              E  d�  dh          E�              -  d�  c�          E�              !  e  c�          E�                e0  bp          F              '  eT  c�          F@              9  ex  dD          Fp              3  e�  c�          F�              ?  e�  d�          F�              ]  e�  e@      �&|�����B��      G               Q  f  e          G0              K  f,  cl          G`              W  fP  d�          G�              i  ft  e�          G�              c  f�  d�          G�              o  f�  ed          H               �  f�  f�          HP              �  g  f<          H�              �  g(  f          H�              {  gL              H�              �  gp  e�          I              �  g�  f�          I@              �  g�  e�          Ip              �  g�  f`          I�  ��D}�;��
S�              �  h   g\          I�              �  h$  g8          J               �  hH  e�          J0              �  hl              J`              �  h�  g�          J�              �  h�  f�          J�              �  h�  g�          J�              5  h�  h|          K                 i   h�          KP              �  iD  hX          K�              �  ih  h4          K�              �  i�  f�          K�              �  i�  h          L              �  i�  h�          L@          �����4;���      �  i�              Lp              �  j  h�          L�                j@  i�          L�                jd  ix          M                 j�  g�          M0                j�  iT          M`              )  j�  i�          M�              #  j�  i0          M�              /  k              M�              e  k<  k          N               M  k`  j�          NP              A  k�  jt          N�              ;  k�  i          N�              G  k�  jP          N�              Y  �W���5|Z|);��  k�  j�          O              S  l  j,          O@              _  l8  j�          Op              }  l\  k�          O�              q  l�  k�          O�              k  l�              P               w  l�  kp          P0              �  l�  l$          P`              �  m  l           P�              �  m4  kL          P�              �  mX  k�          P�              �  m|  l�          Q               �  m�  k(          QP              �  m�              Q�              i  m�  ]�  ��͹$M���{���                         1  n  \�          P              	/  n0              �              		  nT              �                nx              �                n�                            �  n�  ^          @              �  n�  X�          p              =  o  Y�          �              �  o,  n@          �              �  oP  n�                         �  ot  n�          0              J  o�              `              �  o�  Z�          �              T  o�  ^�          ����G���UD�7  �                p  ^�          �              	  p(                             �  pL  b�          P              �  pp  V�          �              �  p�  Z�          �              �  p�  Y          �              �  p�  _�                        �  q   VX          @              (  q$  m�          p              �  qH  p8          �              �  ql  p�          �              �  q�  p�                          �  q�  mD           0              n  q�  \           `      ��W��-�3���          �  q�  q�           �              	B  r   [�           �              $  rD               �              	L  rh  q�          !               	G  r�  q4          !P              	O  r�  X�          !�              �  r�  _�          !�              
)  r�              !�              	�  s  r�          "              	�  s@  Z$          "@              	y  sd  q�          "p              	d  s�  o          "�              	_  s�              "�              	n  s�  ^8          #               ��0Q{T<���Y�  	�  s�  [           #0              	�  t  l�          #`              	�  t<  ^\          #�              	�  t`  \�          #�              	�  t�  ^�          #�              	�  t�  Z�          $               	�  t�              $P              �  t�  m�          $�              �  u              T               	�  u8              $�              	�  u\  p          $�              	�  u�              %              	�  u�  qX          %@              	�  u�  t(          %p              	�  u�  �Ht�Ec�c  o�          %�              
  v  at          %�              
	  v4  n          &               
  vX  ul          &0              �  v|  rx          &`              F  v�  o�          &�              j  v�  [h          Rp              V  v�  ll          R�              `  w              R�              }  w0  r�          S               �  wT  u           S0              O  wx  p�          S`              r  w�              S�              �  w�  ^�          S�              �  w�  r      ���Y��V�dd      S�              
1  x  v�          &�                x,  u�          &�              
<  xP  rT          '               
G  xt  d�          'P              !  x�  WT          '�              '  x�  s�          Q�              /  x�  g�          Q�              7  y  v           R              =  y(  t          R@              �  yL  o`          '�              
O  yp              '�                y�  v�          (              �  y�  st          (@              ?  y�  d           (p  ��җ�K���g��              
W  z   r�          (�                z$              (�              
a  zH  a,          )               �  zl  x�          )0              [  z�  g          )`              4  z�  \@          )�              �  z�              )�              
k  z�  x          )�              �  {   p\          *               
s  {D  w�          *P              
{  {h  [�          *�               e                                                                                                      �8q�_`x��Q                                                                                                                                                                                                                                                                                                                                   e                                          ~�                                                                                                                                                  ����Xo 2���                                                    ~�                                                                                                                                                                                    ~�              *�                               *�                $              +               e                                                                              �$                  �                                                                        V�	r � �*�                                                                          �H                                                                                                                                                      ��                          -  ��              +@              "  �              +p              )  �8              +�                �\              +�               e                                                                                                                  �x�6�S�%2                                                                  �                      �8                          �\                                                                                                                                                                                              S  �(              ,               F  �L              ,0              @  �p              ,`               e                                                                              ��              �h����                      ��                                                              �(                                                      �p                                                                                          ��                                                                  �L                          S  �<              ,�              r  �`              ,�              f  ��              ,�              t  ��              -               x  ��              -P              v  �l�k��T�3  ��              -�               e                                                                                                          ��                                                                      ��                                                                                                                                                                                                                                                  �  ��              -�              S  ��              ��=�'�dPB�  -�               e                                                                                                                                                                              �  ��                                                                              ��                                                                                                              ��                                                  �  ��              .              S  ��              .@              �pW���<��tp  �  ��              .p              �  �              .�               e                                                                                                                                                                                  ��                                                                                                                                                                                                                                              ��  �  ��          �q���d�/"�@      .�              S  �              /                e                                                                                                                                                                                  ��                                                                                                                                                                                                                                              ��  �  ��              /0          �q!�����G��      S  ��              /`               e                                                                                                                                                                                  ��                                                                                                                                                                                                                                                  S  ��              /�               e          �s��Xko���                                                                                                                                                                                                                                          �|                                                                                                                                                                                    ��              /�               e                              ��                              	��@��4�)                                                                                      ��                              �h                                      �H  ��                                                      �l                                              �D                                              ��              �                                 �\              /�              �  ��              0               �  ��              TP              !  ��              0P                ��  
�{|��(c���_&              0�                �              0�                �4              0�              �  �X              1              �  �|              T�               e                                                                                                                                                                                                                                                                                                                  �4                              �s|k�������                                                      �X                              /  �H              1@              6  �l              1p               e                                  ��                                                                  �l          �                                                                       ��                                                      �D                                                                  ��                                          )q���z�'��                                          �h                          g  �8              1�              �  �\              1�              �  ��              2               �  ��              20                ��              2`              m  ��              2�              Q  �  �H          2�              Z  �4  �$          2�              `  �X  ��          3               I  �|              3P               e                                                                                  �� ]�g.��4��                                                                                                                                                                                                                                                                                                                                                                    ���@�� �$                   ����@�����@����@ �(    �                @ �  ֠ � ��   ����� ֠\����@@@@@@@@@@@@@@@@@@@@@@@@@\����@@@@@@@@@@@@@  e�2IR��.rR@@@@@@@@@@@@\��@@@@@@@����`�@@@@@@@@@@@@@@     %�������������   ����                                            �����@������@@@@      0          @����nnnnnnnn����@����������@      �          � � ���@���@Ӊ�����@剅�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@���a���@@@@@@@@@\�   %@    :������������� sd�������� ��  �������������@����@@@    �     �� ������@@@@@@@@@\������@�����@���@����@���������@�����    \������@@@      \�����@@@@      \��@@@@@@@      ����`��         \������@@@      @@@@@@@@@@@@@�@�@Ć��  ���Hrj�=b�^�����M\��]@������M}�����}]@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@@�@�@���������@@M}ǉ������@Ö���������@����@`@����������|�����K��}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@@�@@aa```````````````````````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����  �����(x��p��@@@@@������@@ @@@@@@@@�@@aa@◖��@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@@�@@aa```````````````````````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@@�@���������@@��@@@�@@@@@@@@@@@@@����@@@@������M�������]@������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �������~@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@@�@@aa```````````````````````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@aa@Ô�@ׁ��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@aa```````````````````````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�ŕ���ׁ���@@@@@@@��@@@@@@@@@@@@@@@@@@������M}  R�4�p��"��������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�������@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�������@@@@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�������@@@@@  �˚�T$=w���@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@������@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@���������@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@���������@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@�  �>�"w�E:������@@ @@@@@@@��@�@����������@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�����������@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@����������@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@����������@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  
B��&nx'�S��@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�����������@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@����������@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�������@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@  zM
Z2X c��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�ŕ���ׁ���@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�������@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�������@@@@@@@@@@@@@  �/R�]r޻:Z,@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�������@@@@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@������@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@���������@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@   �e]�/���
�g@@@@@@@��@�@���������@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@����������@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�����������@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@����������@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  K� �vЕ{�77�@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@����������@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�����������@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@����������@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@  �5�͉U�(ԗs�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�������@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@������@@@@@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@\@ؤ�@��@@@@@@@@@@@@@@@@@@@@@  �D7���5�f��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�������@@@@@@@@@@@@@@@@@�@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@\@¨���@י������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�������@@@@@@@@@@@@@@@@@�@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@�  �(Z����V���@@\@¨���@���������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�����@@@@@@@@@@@@@@@@@@@�@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@\@ŧ�������@Ʉ@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@��������@@@@@@@@@@@@@@@��@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��l�O�ny�@@@@������@@@@@������@@ @@@@@@@��@@\@偙����@������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@\@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@���������@@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@\@ؤ�@��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �I���<�W�A�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@������@@@@@@@@@@@@@@@@@@�@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@\@҅�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@���������@@@@@@@@@@@@@@@�@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@\@¨���@י������@@@@@@@@@@@@@@@@@@@@@  ͝�؍�0�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@���������@@@@@@@@@@@@@@@�@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@\@¨���@���������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�������@@@@@@@@@@@@@@@@��@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@\@ŧ�   4���JX��.�n�������@Ʉ@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@����������@@@@@@@@@@@@@��@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@\@م������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@@����������@@@@@@@@@@@@��@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����  !�7ml�UjCtT(��@@@@@������@@ @@@@@@@��@@\@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@��������@@@@@@@@@@@@@@@��@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@\@ֆ����@ŧ�@ā��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@��������@@@@@@@@@@@@@@@��@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  "~`��K��)AS�@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@��������@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@aa@⣙���@����@��ɢ@``````````````````````````````````````````````````K@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@Ĥ�����@@@@@@@@@@@��@@@@@@@@@@@@@��@�@�������M  #<�f�q.�?=E}������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@Ė���@@@@@@@@@@@@@��@@@@@@@@@@@@���@�@�������M}����}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@@@@@@@@@@@@@  $��h���+�p2�@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@�������M\������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@�������M\������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�m�����@@@@@@@@@�@@@@@@@@@@@@@���@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@�  %�y�v�n����"������@@ @@@@@@@��@�@�m������@@@@@@@@�@@@@@@@@@@@@@���@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�m�����@@@@@@@@@�@@@@@@@@@@@@@���@�@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�m��������@@@@@@�@@@@@@@@@@@@@���@�@���M�������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�m�����@@@@@@@@@�@@@@@@@@@@@@@���@�@���M���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  &n��K�7��at�@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@�m�����@@@@@@@@@�@@@@@@@@@@@@@���@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@Ħ����@@@@@@@@@@@@��@@@@@@@@@@@@���@�@�������M}�����}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\@@@�����@@@@@@@@@@@  '4��D<�8E@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@ă����@@@@@@@@@@@@��@@@@@@@@@@@@���@�@�������M}�����}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@aa@@@@@@@@@@@@@@@@@@@  (�f�D�j�]�h@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@Ć�@@@@@@@@@@@@@@@�@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@��@@aa@Ӗ���@����������@``````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@   )Ћ9I�;���@@@@@@@��@�Ⅳ��ׁ��@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�Ù���Ƣ���@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@������@@@@@@@@@@@@@@@@@@@@@@@����@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  *�C��f-`�]�@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�晉��ȅ����@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@㉣��@@@@@@@@@@@@@@@@@@@@@@@@����@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�晉��ׁ���@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  +�h��"���w@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�晉��ׁ���㙅�@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�晉���م�@@@@@@@@��@@@@@@@@@@  ,�/�x�w���c@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�晉��㙁����@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@��  -�jdaD�����#�@�⣁��ׁ��@@@@@@@@��@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ŕ�ׁ��@@@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@⣙���⣁��@@@@@@@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  .��փ�7��'��.@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�晉��ā��@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@¤����@@@@@@@@@@@@@@@@@@@@@@�����@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@Ӆ�@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@  /����;D����n@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�Ó�����Ƣ���@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ɕ�ん�����@@@@@@��@@@@@@@@@@@���@@@@  0�K�b;�aAH@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ǅ�ř�ɕ��@@@@@@@��@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�╄ׇ  1M��u�?Ƙ�Y�Ԣ�@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@����@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@��������@@@@@@@@@@@@@@@@@@@@@@���@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@���Ʉ@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����  2���튾�<�En��@@@@@������@@ @@@@@@���@�@���@@@@@@@@@@@@@@@@@@@@@@@@@@����@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@Ö��������@�����@``````````````````````````````````````````````````@@@@@@@  3>w�\��N��4@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ん�����@@@@@@@@@�@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@ԉ��@���������@````````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@���@@@@@@@@@@@@@@@�@@@@@@@@@@@@@@@@@@@�}��}@@@  4?(J���z=@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@���@偙������@`````````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ׁ��Ֆ@@@@@@@@@@@�@@@@@@@@@@@@@@��@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ׁ��ւ����@@@  5���Ku�8Ї:�@@@@�@@@@@@@@@@@@@@��@�@���M���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@ħւ����@@@@@@@@@@�@@@@@@@@@@@@@@��@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@ħֆ����@@@@@@@@@@�@@@@@@@@@@@@@���@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@ħم�@@@@@@@@@@@@@�@@@@@@@@@@@@@���@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@�  6���}��{z�;������@@ @@@@@@���@�Ӗ�������@@@@@@@@�@@@@@@@@@@@@@���@�@���M����]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ז���≩�@@@@@@@@�@@@@@@@@@@@@@@��@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�兙�◁��@@@@@@@@�@@@@@@@@@@@@@@��@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  7��3��s��U�@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�Ö��@@@@@@@@@@@@@�@@@@@@@@@@@@@@��@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�Ӆ��ԁ����@@@@@@@�@@@@@@@@@@@@@@��@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�㖗ԁ����@@@@@@@@�@@@@@@@@@@@@@@��@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  8r�/���z�B�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ׁ��扄��@@@@@@@@�@@@@@@@@@@@@@@��@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ׁ��ȅ����@@@@@@@�@@@@@@@@@@@@@@��@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@  92�i�D��?�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ą�����Ɩ��@@@@@@�@@@@@@@@@@@@@@@@@@@}Ö�����}@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�Ɩ��@@@@@@@@@@@@@�@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@   :)K^.���d��@@@@@@���@@aa@י�����@������@````````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ׇ�⣢@@@@@@@@@@���@@@@@@@@@@@@@@@@@@Ֆ֗�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@і�Ղ�@@@@@@@@@@@@@@@@@@@@@@@@@��@@@֥�����Mׇ�⣢z���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ;���Vh�yRh@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  <L,�/#S��=�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@Ⅳ��@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���~����������@@@@@@@@@@@@@@@@@@@@  =6ITX�YW�esH@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������@@ @@@@@@���~�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�@@@@�@@@@�@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������@@ @@@@@@���~�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�@@@@�@@���@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������@@ @@@@@@���@@@Ⅳ��ׁ��@M]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@��  >zaCe�p,�h���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@Ù����@���@���@������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@Ù���Ƣ���@M������]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ?���0s��Ђ&� @@@@������@@@@@������@@ @@@@@@���@@@aa@ɕ��������@����������@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@ん�����@~@ɕ�ん�����M]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@晉��@��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  @jY�y��F�[�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ȅ����M�����]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ׁ���M]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ׁ���㙅�M]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉���م�M]^@@@@@@@@@@@@@@@@@@@@@@@@  A��9 k��4��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��㙁����M]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@�����@������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@Ó��  B�5�A�r�������Ƣ���@M]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@\����@~@\��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����  C�k �}��[��@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@  D�$� �&�9�E4@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@Ⅳ@ׁ��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�Ⅳ��ׁ��@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�Ⅳ��ׁ��@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@  Eh���� �@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@��@���������@~@}\����}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@������^@@@  F�4'�قV���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@����@�������@L~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@���������@~@}\����������}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@����@�������@L~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@�  G|����U���9������@@ @@@@@@���@@@@@@@@@���������@~@}\������������}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@���������@~@}\������������}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  HT����K�7j�@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@����@���������@~@}\����������}^@@@@@@@@@@@@@@@@@@@  Ii�����Or�G@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@ׁ��扄��@@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@ׁ��ȅ����@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@ז���≩�@@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@兙�◁��@@~@��^  J��#t����
^�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@Ö��@@@@@@@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@Ӆ��ԁ����@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@㖗ԁ����@@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@   K>��X�gĐ��@@@@@@���@@@@@����@���������@~@}\�����������}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@ׁ��扄��@@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@ׁ��ȅ����@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@ז���≩�@@~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  L���Oh2�F�<@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@兙�◁��@@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@Ö��@@@@@@@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@Ӆ��ԁ����@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@㖗ԁ����@@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  MŚYfc���"�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@����@���������@~@}\������������}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@ׁ��扄��@@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@ׁ��ȅ����@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@ז���≩�@@~@��^@@@@@@@@  N򁲈C�7Q���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@兙�◁��@@~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@Ö��@@@@@@@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@Ӆ��ԁ����@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@��  O�Y�R��Yq�O�@@@@@@@㖗ԁ����@@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@����@���������@~@}\������������}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@ׁ��扄��@@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@ׁ��ȅ����@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@  P�ī���m#I�:@@@@������@@@@@������@@ @@@@@@���@@@@@@@ז���≩�@@~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@兙�◁��@@~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@Ö��@@@@@@@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@Ӆ��ԁ����@~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  Q��JDC];���@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@㖗ԁ����@@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@����@���������@~@}\������}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@ׁ��扄��@@~@����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@ׁ��ȅ����@~@�����������^@@@@@@@  R��t	���g@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@ז���≩�@@~@����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@兙�◁��@@~@����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@��@�Ö��@~@`�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@  S�瓰3uY��ͬ�@@Ö��@~@�������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@Ö��@@@@@~@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@����  T[�C�"1=k���@@@@@������@@ @@@@@@���@@@@@@@Ӆ��ԁ����@~@�����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@㖗ԁ����@@~@����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  U��=Ґu��d��@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@��@�֙����@~@}\���������}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@ׁ��扄��@@~@�ׁ��ȅ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@ׁ��ȅ����@~@�ׁ��扄��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  VB��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�Ⅳ��ׁ��@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@  W������X�S>��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@Ù����@��@�����@���@������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@�  Xv��ɭ���-������@@ @@@@@@���@�Ù���Ƣ���@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�Ù���Ƣ���@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@������@@@@@@@@@@@@@@@@@@@@@@@����@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  Y��x�ʨ��%(�@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�Ɖ��Ձ��@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ř�Ԣ�@@@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  Z�'��Ԝ�ް@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@Ɖ��Ձ��@~@l����M������]@N@�}��}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@È���@�������@���  [��ۃD�(s�JN���@����@������@��@���K@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@��@~@����Ml����MƉ��Ձ��]@z@�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@Ɇ@⣙���@����@������k@����@������@���@������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@   \�C���{�'�,,@@@@@@���@@@Ɇ@��@Ln@`�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@Ɇ@�����M��]@~@`�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@ř�Ԣ�@~@}�����M]@������K@}@N@����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@ŕ�Ɇ^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ]����8���E�Q�@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@Ɇ@������Ml����MƉ������]]@~@`�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@ř�Ԣ�@~@}������M]@������K@}@N@����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@ŕ���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@ŕ�Ɇ^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ^:ꢕu�sZN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@��@������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@��@ř�Ԣ�@Ln@}@}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@╄ׇ�Ԣ�@M}\������}z}Ù��  _�G�E�Uh�����Ƣ���}z@}@}@z@ř�Ԣ�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@ŕ���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@֗��MÙ����]@������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@��  `��2�k���@@@��@~@����Ml����MƉ������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@z@�m�����@N@�m������@N@�m�����@N@�m��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@z@�m�����@N@�m�����@z@���]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@Ɇ@��@~@`�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@  a�i��&=r^C��c@@@@������@@@@@������@@ @@@@@@���@@@@@ř�Ԣ�@~@}����M]@������K@}@N@����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@ŕ�Ɇ^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@��@������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  b��Saoh�\�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@��@ř�Ԣ�@Ln@}@}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@╄ׇ�Ԣ�@M}\������}z}Ù���Ƣ���}z@}@}@z@ř�Ԣ�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@ŕ���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  c�|c0y�2ɨ�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�Ù���Ƣ���@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@  d��C<���"@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@晉��@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����  eX���n�XXZG���@@@@@������@@ @@@@@@���@�晉��ā��@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�晉��ā��@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@¤����@@@@@@@@@@@@@@@@@@@@@@�����@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@Ӆ�@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  fq�{�X���78@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@������@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@ħ�����@@@@@@@@@@@��@@@@@@@@@@@@@@@@@@�������M}m������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\@@@�����@@@  g�������b5�)�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�¨����@@@@@@@  h��h���q���d@@@@�@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ř�Ԣ�@@@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@�  i�;�6��P@R"������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@�������@��@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@������@Ml����M¤����]zl����Mん�����]zӅ�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  j&����TP����@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@�����@����@��@������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@¨����@~@�����M��zl����M¤����]zӅ�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@Ɇ@¨����@Ln@Ӆ�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@ř�Ԣ�@~@}�����M]@������K@}@N@����������^@@@@@@@@@  k��>�V��9	�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@ŕ���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@��������@�����@��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@�ֆ����@N~@¨����^@@  l�P�Q��(�]��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@   mq+ }Ĭ����@@@@@@���@�晉��ā��@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@晉��@������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  n��k��/|��je@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�晉��ȅ����@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�晉��ȅ����@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@㉣��@@@@@@@@@@@@@@@@@@@@@@@@����@@@�����@@@@@@@@@@@@@@@@@@@  o]�פ^�w���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@Ù������ā��@@@@�@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@œ�����@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  pUǛ�I/��j���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@�������@���@�������@���@����@ȉ�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@��  qYݭk ��m��Ci�@@@晉��ā��M}l���`�K�}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}l}@N@�}��������}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@��������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  r2�(ƃ�{��@@@@������@@@@@������@@ @@@@@@���@@@Ӗ�������M�]@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}�@�@���}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}LL}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@Ù������ā��@~@l����Ml����M]z\����]Nl����Ml����M]z\����]^@@@@@@@@@@@  s��cW��z%�u:�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}aÙ������ā��@M�z}@N@Ù������ā��@N@}]}N@��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}aי������@M�������@��K�@M����@���Ö���k@����]]}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@œ�����@~@}a㉣��@M}@N@l����M㉣��]@N@}]}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��Mœ�����zl���Ml�����Mœ����  t�w�#5rs]��`�]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}nn}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}������}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@�  u=�Ǝ�}��9o���@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@Ӗ�������M�]@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}�@�@���}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}LL}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����  v�tjLN"vs�����@@@@@������@@ @@@@@@���@@@晉��ā��M}a㨗�@aÁ�����}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}aׁ���@�@�@�}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}nn}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}������}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  wn�A]y�C磻�@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@Ӗ�������M�]@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}�@�@���}N��z�]^@@@@@@@@@@@@@@@@@@  x1�I'!�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}LL}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}a㨗�@aƖ��}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}a⤂����@a㨗��}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}a  yt��s�P�5Ձ��@a��}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@��@���������@~@}\���}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@Ɩ��@~@ą�����Ɩ��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@�  z�.�T,��������@@ @@@@@@���@@@@@Ɩ��@~@���������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@œ�����@~@}a��Ɩ��@a}@N@l����MƖ��]@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  {PPr_�#���|@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}aŕ������@a払����ŕ������}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}nn}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}������}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  |?�K�RG�k1I,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@����@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@Ӗ�������M�]@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}�@�@���}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}LL}N��z�]  }�<��\!S%�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}@@aƖ��@LL@a��@�@�@�@nn}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}@@aי��Ⅳ@�@a���@aㅧ�@�}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}nn}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@   ~�x��B{��a�@@@@@@���@@@晉��ā��M}������}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�晉��ȅ����@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��I:�Ȁ����@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@晉��@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN  ��V�MQ\�z'�NNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�晉��ׁ���@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�晉��ׁ���@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@œ�����@@@@@@@@@�@@@@@@@@@@@  �"	�Ϻ!V��T@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@���⣙���@@@@@�@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@��  ��?��[�KA���S�@�@�@@@@@@@@@@@@@@@�@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@�@@@@@@@@@@@@@@@�@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@�@@@@@@@@@@@@@@@�@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@ׁ���������@@@@@�@@@@@@@@@@@@@@@@@@@}�M]}@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �7��_�Ĳ���@@@@������@@@@@������@@ @@@@@@���@�@ׄ�ㅧ�@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �/�h~Vz��LX\@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@����@��������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@���@���@l���M��������]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@aa@����@�@���@����@@@@@@@@@@@@@@@@  �b�0W�m�jT-8@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@�����������@~@⣁��ׁ��M]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@aa@����@�@�����@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@����@��������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@��  �4����q0dOտ�@���@l���M��������]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@晉��ā��M}M}z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@ׄ�ㅧ�@~@����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@aa@������@�����������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����  ��8dx`D�/�,���@@@@@������@@ @@@@@@���@@@@@@@���@�@~@�@��@l���Mׁ���������]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@�@~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@�@~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@���@�@~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ����@��*���@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@�@~@l����Ml�����Mׁ���������z�z�]zl�����Mׄ�ㅧ�z�N�]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@��@�@n@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@�@N~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@ׄ�ㅧ�@~@l�������M}�}zׄ�ㅧ�z�z�  ��"
e�C_����]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@�@N~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@������^@  ��Y�lj��N>@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@aa@�����@�����@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@晉��ā��Ml�����Mׄ�ㅧ�]zl���Ml�����Mׄ�ㅧ�]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@晉��ā��M}]}}}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@�  ���-�g�'��M�����@@ @@@@@@���@@@@@@@aa@����@����@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@����@��������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@��@���@l���M��������]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@aa@������@����@�����������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �{܏�j�9U<�E@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@����@����@~@}�}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@ŕ�ׁ��M�����������]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@�����������@~@⣁��ׁ��M]^@@@@@@@@@@@@@@@@  ����?|���T��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@����@����@~@}�}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@晉��ā��M}M]}}}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@����@����@~@}`}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@晉��ā��M}  ����(��8�;�RM]}}}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@晉��ā��M}M]}}}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@   ��k����F9+@@@@@@���@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@aa@�����@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@ŕ�ׁ��M�����������]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��,�^O��Uj�@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@�����@��������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��Ei��P����n@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�晉��ׁ���@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@⣁��@����@@@@@@@@@@@@@@@@  �eS>��'��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�⣁��ׁ��@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�⣁��ׁ��@@@@@@@@��@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@��  ��di���6��6�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@����ז�@@@@@@@@@�@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@œ�����@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��ٱ��2�H�R@@@@������@@@@@������@@ @@@@@@���@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@�ւ����@N~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �7���e��m�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@Ӗ�������M�ւ����]@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@����Ֆ@N~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@ׁ��ւ����M����Ֆ]@~@�ւ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@œ�����@~@l����M�ւ����]@N@}@�@���}@  ����\��a}Q�N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}LL}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}a㨗�@aׁ��}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉�  �����\˗�E��ā��M}aׁ����@�@�@�}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}aم�������@�@�@�}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@�ւ����@N~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@œ�����@~@}aÖ������@}@N@l����M�ւ����]@N@}@�@�}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����  ����D�������@@@@@������@@ @@@@@@���@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}nn}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}������}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �`�"0��|��]��@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@Ӗ�������M�ւ����]@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@œ�����@~@l����M�ւ����]@N@}@�@���}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��
�B�<���Ն@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}LL}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@œ�����@~@}aӅ����@}@N@l����M�ւ����@N@�]@N@}@�@�}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@  ����R��p��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}nn}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}������}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@����ז�@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@�  ��84�_D�_��������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@��@�����@�@����@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}��}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �"�����qez@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@���@�������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@œ�����@~@}a��@}@N@l����M�����≩�]@N@}@�}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �1������k��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@���@�������@M�k�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@œ�����@~@}�@�@�@�@}@N@l����M����ԁ����]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@}@}@N@l����M����ȅ����@`@���ԁ����]@N@}@�}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��Mœ�����zl�  �}����>�u1M��Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@���@��������@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@œ�����@~@l����M����◁��]@N@}@��}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@   ��6�߾Q�C��@@@@@@���@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@������@����ז�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��C�!��F[�@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�⣁��ׁ��@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN  ����&�]�W�u	NNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@ŕ�@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ŕ�ׁ��@@@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ŕ�ׁ��@@@@@@@@@@��@@@@@@@@@@  ��
&���P�nN�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@⣙���⣁��@@@@@@@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@œ�����@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@��  ���vt:������ �@�@⣙���ŕ�@@@@@@@�@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@aa@��@����@���@����@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ���P. ��^m0�@@@@������@@@@@������@@ @@@@@@���@@@@@晉��ā��M}��}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@������ŕ�@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@晉��ā��M}���������}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@晉��ā��M}������}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �&D���)e�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@�ւ����@N~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@Ӗ�������M�ւ����]@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ���wɋt�_��%@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@œ�����@~@l����M�ւ����]@N@}@�@���}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@œ  ��)zl~���\Lۅ����@~@l����M⣙���ŕ�@`@������⣁��]@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@晉��ā��M}������}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����  ��	��ԥ�[.��@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ŕ�ׁ��@@@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �������RE�@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@晉��@�����@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�晉��ׁ���㙅�@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@  �5s<exDY�'�=@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�晉��ׁ���㙅�@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@�@@@@@@@@@@@@@@@�@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@  ��kpv-�?ى�|Q@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@œ�����@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@�  ��;�6#u�/��(�����@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@Ӗ�������M�]@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}�@�@���}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}LL}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �+�`�����@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}a㨗�@aׁ���}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@������@����@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@œ�����@~@}aÖ���@}@N@l����M����Ֆ]@N@��^@@@@@@@@@@@  �x���!q�D��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@������@���������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@œ�����@~@}aԅ����  ���I^<����@�@�@�@}@N@l����M����扄��]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@}@}@N@l����M����ȅ����]@N@}@�}@N��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@   �0��r�j��^@@@@@@���@@@aa@������@������@���������@��@����@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}a҉��@�}z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@���@�@~@�@��@����Ֆ^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@��@l���M�z��]@~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��l�a�M� �2�@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@晉��ā��M��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@œ�����@~@}@}@N@l����Mׁ��ւ����M�]]@N@}@�@�}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@  �q@�0(�m��W@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}@�}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}nn}N��z�]^@@@@@@@  �����+	�|L@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}������}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@��  ���1?���yA�!��@�晉��ׁ���㙅�@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@晉��@�م�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �?�J`��u��t��@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�晉���م�@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�晉���م�@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��r}��X��G'@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@�@@@@@@@@@@@@@@@�@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@œ�����@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��K��
���.�(@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@�����@�م�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@�م�  �ʙgӀD����
@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}����}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@KKK@������@��@�������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����  ��Ys��iUe^����@@@@@������@@ @@@@@@���@@@œ�����@~@}�@}@N@l����M�ւ����@N@�]@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@KKK@����@�����@`@����@��@������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ���R��k��p��@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@œ�����@~@}����������@�����@�@}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@KKK@�م�@�������@@@@@@@@@@@@@@@@@@@@@@@@@  �Op� e*��7A@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@���@�@~@�@��@�ւ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@œ�����@~@l����Ml�����Ml���MӖ�������M�]z��z�]z}�}]]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@}@�����@�@}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@晉��ā��M  ��6	�:\�庙œ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@�  ��9f#?�w�k�gp�����@@ @@@@@@���@�晉���م�@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@晉��@�������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �	��!��σ�k�;@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�晉��㙁����@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�晉��㙁����@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �z�-�Pv�Om&mP@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@œ�����@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@  ���?h���]⋘@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}�������}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}LL}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@   �1��,!�pa�@@@@@@���@@@aa@�����@������@��@�������@��@�م�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@œ�����@~@}a≩�@}@N@l����M�ւ����@N@�]@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}aٖ��@�@�@�}N��z��]^@@@@@aa@���������@��@Á�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��nq_�w5�K)8@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}aɕ��@�@�@�}N��z��]^@@@@@aa@���������@��@ɕ��@����������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}nn}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@������@��@�م�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �+� Y䆖q�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}���������}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@œ�����@~@l����M�م�]@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ������.h��_VI@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@aa@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@晉��ā��M}ll���}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@��  ��t������@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�晉��㙁����@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  Ǉ���x���F@@@@������@@@@@������@@ @@@@@@���@@aa@Ó���@���@������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�Ó�����Ƣ���@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�Ó�����Ƣ���@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �.��ܧ�Ț�`n@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ř�Ԣ�@@@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@Ɇ@�����M��]@~@`�^@@@@@@@@@@@@@@@@@@  � ���n�=Ώ`@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@ř�Ԣ�@~@}�����M]@������K@}@N@����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@╄ׇ�Ԣ�@M}\������}z}Ó���Ƣ���}z@}@}@z@ř�Ԣ�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@ŕ�Ɇ^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@a���`  �/vr��(l['_�Z����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�Ó�����Ƣ���@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����  ˉe@/���H�h���@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@ɕ��������@あ��@ł����@`n@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ɕ�ん�����@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �|`�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ɕ�ん�����@@@@@@��@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@Ö�����@�@Ǚ�����@È�������@⣙���@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@��������@@@@@@@@@@��@@@@@@@@@@@@@@@@@@������M}  ͏�X<�*\7�����������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@������@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@���@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@��@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@��@@@@@@@@@@  ���]�,o�B�@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@������@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@���@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@������@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@�  Ϸl�ȹ�b�a��������@@ @@@@@@���@�@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@��@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ���q��t�X��H@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@���������@@@@@@@@@��@@@@@@@@@@@@@@@@@@������M}��������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@��������@@@@@@@@@@@@@@@@@@@@����@@@@�������M\�������  �Y ih}�O��g]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@����¨���@@@@@@@@@@@@@@@@@@@@@@��@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@����Ɩ����@@@@@@@@@@@@@@@@@@@@��@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@����і�Ձ��@@@@@@@@@@@@@@@@@@@��@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@����і�ɕ�@@@@@@@@@@  �"P��b�P�@@@@@@@@@@��@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@���ř���@@@@@@@@@@@@@@@@@@@@@���@@@@�������M\�������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@��������@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@@�����@@@@@@@@@@@@@@@@@@@@@@@@@��@�@�������M��������z���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@   ��C=���xL �:�@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@����������@������@���@�������@���@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ん�����@@@@@@@@@�@@@@@@@@@@@@���@@@@���M\����}��}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�んł����@@@@@@@@�@@@@@@@@@@@@���@@@@���M\����}��}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  Զ�o2g0fF�k@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@���@@@@@@@@@@@@@@@�@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@���@@@@@@@@@@@@@@@�@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@���@@@@@@@@@@@@@@@�@@@@@@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ����*��܂�*"@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@����������@������@`@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@��偓��@@@@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@�偓��@@@@@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ։�5�݈:��~�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@aa@���@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@��������@M��������zl���M��������]z}��������}z}\}z}@}z�����]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@��  ו��-ٯ[@�ZD�@@@@aa@������@�@����������@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@���@�偓��@~@�@��@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@l�����Mんł����z�偓��N�z�]@~@�偓��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@  �z�w���+��7j@@@@������@@@@@������@@ @@@@@@���@@@@aa@������@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@�������@M�����z�zんł����z���z���z�z�z���zん�����z��z��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@aa@������@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@������@ん�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ���L5�7���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�ɕ�ん�����@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ڈK��׹eև(@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@ǅ�@�@�����@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@ׇ����  �z�<Y�8t��n�����@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@ć���������@@@@@@@��@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@ć�������@@@@@@@@@��@@@@@@@@@@@@@@\@@@�������M}mm�����}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@Ģ�������@@@@@@@@@��@@@@@@@@@@@@@@\@@@�������M}��������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����  ܈�Sc1�.�O�n��@@@@@������@@ @@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@ą�����@@@@@@@@@@@�@@@@@@@@@@@@@���@�@�����M������m�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@������m�@~@��������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ���wÒ��ǩ�@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@م����@l����Ml�����M������@z@}�}]]@N@}@z@}@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@l���M��������M������]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@ׇ���������@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@  ޙ}0x(��C�YE@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aa@⅕�@י�����@ԅ�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@aaNNNNNNNNNNN  �u�}�)��>NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�╄ׇ�Ԣ�@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�╄ׇ�Ԣ�@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@���㨗�@@@@@@@@@@@@@@@@@@@@@@@���@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@�  ��\��0���I�����@@ @@@@@@���@�@��������@@@@@@@@@@@@@@@@@@@@@@���@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@���Ʉ@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@���ř�@@@@@@@@@@@@@@@@@@@@@@@����@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��L�dt\�K!�@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@��������@@@@@@@@��@@@@@@@@@@@@@@@@@@������M}��������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@@ԅ�����Ʉ@@@@@@@@@@@@@@@@@@@@@�@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@@ԅ�����Ɖ��@@@@@@@@@@@@@@@@@@��@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@@ԅ�����ā��@@@@@@@@@@@@@@@@@���@@@@�����@�������M\�  �Z��V���F4ہ�����]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@@ԅ�����ā���@@@@@@@@@@@@@@@@@@��@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@@ԅ�����㨗�@@@@@@@@@@@@@@@@@@��@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@@Á��⣒ŕ���@@@@@@@@@@@@@@@@���@@@@�����@�������M\�������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@@Á��⣒Ö���@@@@@@@  �~�6�{q���@@@@@@@@@@@��@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@@ԅ�����҅�@@@@@@@@@@@@@@@@@@@@�@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@@���ř���@@@@@@@@@@@@@@@@@@@@���@@@@�������M\�������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@   �%$������ԤR@@@@@@���@�@��Ԣ�@@@@@@@@@@@�@@@@@@@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�@���Ԣ�@@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��;U��ZUJD�T@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@��@���Ʉ@Ln@}@}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@��Ԣ�@@~@���Ʉ^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@���Ԣ�@~@���ř�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ���5�#[��Q�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@��@���㨗�@~@}\������}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@��Ԣ�@@~@}�������}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@���Ԣ�@~@}ř���@}@N@l���  �'J����F4������M��������]@N@}@z@}@N@���ř�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@���Ԣ�@~@���ř�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@������@@@@@������@@ @@@@@@���@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@��  ���3X��SO�U��@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@��������@M��Ԣ�z@}�������@@@����}@z@���Ԣ�@z@l���M���Ԣ�]@z@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@���㨗�@z@}\������}@z@�@z@}@}@z@�����]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �p=��AX�Vl��@@@@������@@@@@������@@ @@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@���@�╄ׇ�Ԣ�@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������@@@@@������@@ @@@@@@@@@\����@���������@����      m����m����m���  m����m����m���  �����@@@@@     ꂯ5�$��ھ��   @@@@@@          �#:��CK        ������@@@@      \����nnnnnnnn����@����������@        :    � ����  @       �    �  (  �  8  �  H  �  X  �  h  �  	x  
   
�    �     �  0  �  @  �  P  �  `  �  p  �  �    �    �  (  �  8  �  H  �  X  �  h  �  x     �    �     �  0  �  @  �   P   �  !`  !�  "p  "�  #�  $  $�  %  %�  &(  &�  '8  '�  (H  (�  )X  )�  *h  *�  +x  ,   ,�  -  -�  .   .�  /0  /�  0@  0�  1P  1�  2`  2�  3p  3�  4�  5  5�  6  6�  �#'m��!���  7(  7�  88  8�  9H  9�  :X  :�  ;h  ;�  <x  =   =�  >  >�  ?   ?�  @0  @�  A@  A�  BP  B�  C`  C�  Dp  D�  E�  F  F�  G  G�  H(  H�  I8  I�  JH  J�  KX  K�  Lh  L�  Mx  N   N�  O  O�  P   P�  Q0  Q�  R@  R�  SP  S�  T`  T�  Up  U�  V�  W  W�  X  X�  Y(  Y�  Z8  Z�  [H  [�  \X  \�  ]h  ]�  ^x  _   _�  `  `�  a   a�  b0  b�  c@  c�  dP  d�  e`  e�  fp  f�  g�  h  h�  i  i�  j(  j�  k8  k�  lH  l�  mX  m�  nh  n�  ox  p   p�  q  q�  r   r�  s0  s�  t@  t�  uP  u�  v`  v�  wp  w�  x�  y  y�  z  z�  �2ǖ\����w��  {(  {�  |8  |�  }H  }�  ~X  ~�  h  �  �x  �   ��  �  ��  �   ��  �0  ��  �@  ��  �P  ��  �`  ��  �p  ��  ��  �  ��  �  ��  �(  ��  �8  ��  �H  ��  �X  ��  �h  ��  �x  �   ��  �  ��  �   ��  �0  ��  �@  ��  �P  ��  �`  ��  �p  ��  ��  �  ��  �  ��  �(  ��  �8  ��  �H  ��  �X  ��  �h  ��  �x  �   ��  �  ��  �   ��  �0  ��  �@  ��  �P  ��  �`  ��  �p  ��  ��  �  ��  �  ��  �(  ��  �8  ��  �H  ��  �X  ��  �h  ��  �x  �   ��  �  ��  �   ��  �0  ��  �@  ��  �P  ��  �`  ��  �p  ��  ��  �  ��  �  ��  홊��k�@s�>  �(  ��  �8  ��  �H  ��  �X  ��  �h  ��  �x  �   ň  �  Ƙ  �   Ǩ  �0  ȸ  �@  ��  �P  ��  �`  ��  �p  ��  ̀  �  ΐ  �  Ϡ  �(  а  �8  ��  �H  ��  �X  ��  �h  ��  �x  �   ֈ  �  ט  �   ب  �0  ٸ  �@  ��  �P  ��  �`  ��  �p  ��  ހ  �  ߐ  �  �  �(  �  �8  ��  �H  ��  �X  ��  �h  ��  �x  �   �  �  �  �   �  �0  �  �@  ��  �P  ��  �`  ��  �p  ��  �  �  �  �  �  �(  �  �8  ��  �H  ��  �X  ��  �h  ��  �x  �   ��  �  ��  �   ��  �0  ��  �@  ��  �P  ��  �`  ��  �p  ��  �  �  �  ��M�g�Z��ճo� ( � 8 � H � X � h � x 	  	� 
 
�   � 0 � @ � P � ` � p � �  �  � ( � 8 � H � X � h � x   �  �   � 0 � @ � P �  `  � !p !� "� # #� $ $� %( %� &8 &� 'H '� (X (� )h )� *x +  +� , ,� -  -� .0 .� /@ /� 0P 0� 1` 1� 2p 2� 3� 4 4� 5 5� 6( 6� 78 7� 8H 8� 9X 9� :h :� ;x <  <� = =� >  >� ?0 ?� @@ @� AP A� B` B� Cp C� D� E E� F F�  �0��5�4I2� G( G� H8 H� IH I� JX J� Kh K� Lx M  M� N N� O  O� P0 P� Q@ Q� RP R� S` S� Tp T� U� V V� W W� X( X� Y8 Y� ZH Z� [X [� \h \� ]x ^  ^� _ _� `  `� a0 a� b@ b� cP c� d` d� ep e� f� g g� h h� i( i� j8 j� kH k� lX l� mh m� nx o  o� p p� q  q� r0 r� s@ s� tP t� u` u� vp v� w� x x� y y� z( z� {8 {� |H |� }X }� ~h ~� x �  �� � �� �  �� �0 �� �@ �� �P �� �` �� �p �� �� � �� � ��  ����ڃ㛋��� �( �� �8 �� �H �� �X �� �h �� �x �  �� � �� �  �� �0 �� �@ �� �P �� �` �� �p �� �� � �� � �� �( �� �8 �� �H �� �X �� �h �� �x �  �� � �� �  �� �0 �� �@ �� �P �� �` �� �p �� �� � �� � �� �( �� �8 �� �H �� �X �� �h �� �x �  �� � �� �  �� �0 �� �@ �� �Pnnnnnnnn����@����������@      �         Ơ�������@⣁������@剅�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����`�@@@@@@@@@@@@@@\�   %@   Q������������� sd�������� Ơ��������  ������^�!�4�����@����������@ �     Q    ֠���� � ��  v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �  �N�ifoxC㋾      v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v   �     v        v       v       v       v       v       v       v       v       v  	     v  
     v       v       v       -       -       -        -  #     -  $     -  %     -  &     -  '     -  (     -  )     -  *     -  -     -  �	-����I����  .   
  -  /     -  2     -  5     -  6     -  7     -  :     -  ;   
  -  <     -  @     �  E     �  V   
  �  Y     �  Z     �  [     �  \     �  _     �  c     �  h     �  r   
  �  s   
  �  v     �  w   
  �  x   
  �  y     �  z   
  �  {   
  �  |     �  }   
  �  ~   
  �     
  �  �     �  �   
  �  �   
  �  �   
  �  �   
  �  �   
  �  �   
  �  �     �  �   
  �  �   
  �  �   
  �  �   
  �p�Tjxh���  �  �   
  �  �     �  �     �  �     �  �     �  �     �  �     �  �     �  �   
  �  �   
  �  �   
  �  �   
  �  �     �  �   
  �  �   
  �  �   
  �  �   
  �  �   
  �  �   
  �  �     �  �     �  �     �  �     �  �     �  �     �  �     �  �   
  �  �     �  �     �  �     �  �     �  �     �  �     �  �     �  �     �  �     �  �     �  �     �  �     �  �     �  �     �  �     �  �  �r9�,��m�X     �  �   
  �  �   
  �  �     �  �     �  �     �  �     �  �   
  �  �     �  �     �  �     �  �   
  �  �     �  �     �  �   
  �  �   
  �  �     �  �     �  �     �  �     �  �   
  �  �     �  �     �  �     �  �     x  �     x  �     x  �     x  �     x  �     x  �     x  �   
  x  �   
  x      
  x     
  x     
  x       x       x     
  x     
  x     
  x  	     x  
     x  ��ð��Ng�B     
  x     
  x       x     
  x     
  x     
  x       x     
  x       x     
  x       x     
  x  "     x  #   
  x  %     x  (     5  -     5  6   
  5  7     5  8   
  5  9   
  5  ;     5  <     5  >     5  ?   
  5  A     5  B   
  5  D   
  5  G     �  L     �  U     �  V   
  �  W   
  �  X   
  �  [     �  \   
  �  _     �  a   
  �  d   
  �  e     �  f     �  g   
  �  h     ���Ξ���
jN%  �  i     �  j   
  �  k     �  k     �  m   
  �  n   
  �  o   
  �  r     �  w     �  �     �  �   
  �  �     �  �   
  �  �     �  �   
  �  �     �  �     �  �   
  �  �     �  �     �  �     �  �     �  �   
  �  �   
  �  �     �  �   
  �  �   
  �  �   
  �  �   
  �  �   
  �  �     �  �   
  �  �   
  �  �     *  �     *  �     *  �     *  �   
  *  �     *  �     H  �     H  �   
  H  �  ��f��.�(�p&     H  �     H  �     H  �     H  �   
  H  �     H  �     C       C       C  	     C       w       w  (     w  )     w  *     w  +     w  +     w  ,     w  -     w  .     w  /     w  /     w  0     w  1     w  2     w  4   
  w  8       BA         �         �         �         �   
      �   
      �         �   
      �   
      �   
      �   
      �   
      �   
      �         �       BB   nnnn  ��P�J��[+����@����������@@      �       �P �P@@@ � ����         F      \      d      �      �      �      �        	     
       %     .     2     B   nnnn���@����������@@     
�  Q    � �@@@  @ �      B  �   C  �   D  �   E  �   F  �   G  �   H  �   I  �   J  �   K  �   L  �   M  �   N  �   O  �   P  �      �      �      �      �      �      �      �      �    	  �    
  �      �      �      �      �      �      �      �      �      �      �   �7���.��/�     �      �      �      �      �      �      �      �      �      �      �       �    !  �    "  �    #  �    $  �    %  �    &  �    '  �    (  �    )  �    *  �    +  �    ,  �    -  �    .  �    /  �    0  �    1  �    2  �    3  �    4  �    5  �    6      7     8     9     :     ;     <     =     >     ?     @ 
    A     B     C     D     E     F     G !    H $    I %    J &    K '    L (    M )    N *    O +    P .    Q /    R 0    S 3    T 6   ����:q�/_y�|l   U 7    V 8    W ;    X <    Y =    Z A    [ F    \ W    ] Z    ^ [    _ \    ` ]    a `    b d    c i    d s    e t    f w    g x    h y    i z    j {    k |    l }    m ~    n     o �    p �    q �    r �    s �    t �    u �    v �    w �    x �    y �    z �    { �    | �    } �    ~ �     �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �   �Gs r��D��~�   � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    �      �     �     �     �     �     �     �     �     � 
    �     �     �     �     �    ��A�Ap~N;Ԯ�   �     �     �     �     �     �     �     �      � #    � $    � &    � )    � .    � 7    � 8    � 9    � :    � <    � =    � ?    � @    � B    � C    � E    � H    � M    � V    � W    � X    � Y    � \    � ]    � `    � b    � e    � f    � g    � h    � i    � j    � k    � l    � l     n    o    p    s    x    �    �    �    �   	 �   
 �    �    �    �    �    �    �    �    �    �    �   �r�<f��q�=�   �    �    �    �    �    �    �    �    �    �    �     �   ! �   " �   # �   $ �   % �   & �   ' �   ( �   ) �   * �   + �   , �   -    . 	   / 
   0    1    2 )   3 *   4 +   5 ,   6 ,   7 -   8 .   9 /   : 0   ; 0   < 1   = 2   > 3   ? 5   @ 9   A :   Qnnnn���@����������@@     
�  Q    ������@@@  @ �   �      �      �      �      �      �      �      �      �    	  �    
  �      �   ���,H��n�ج�     �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �       �    !  �    "  �    #  �    $  �    %  �    &  �    '  �    (  �    )  �    *  �    +  �    ,  �    -  �    .  �    /  �    0  �    1  �    2  �    3  �    4  �    5  �    6      7     8     9     :     ;     <     =     >     ?     @ 
    A     B     C     D     E     F     G !    H $    I %    J &    K '    ���2�P�C��   L (    M )    N *    O +    P .    Q /    R 0    S 3    T 6    U 7    V 8    W ;    X <    Y =    Z A    [ F    \ W    ] Z    ^ [    _ \    ` ]    a `    b d    c i    d s    e t    f w    g x    h y    i z    j {    k |    l }    m ~    n     o �    p �    q �    r �    s �    t �    u �    v �    w �    x �    y �    z �    { �    | �    } �    ~ �     �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �   7��s�y�����   � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    �      �     �     �     �     �    ��X$.�Dڀ   �     �     �     � 
    �     �     �     �     �     �     �     �     �     �     �     �     �      � #    � $    � &    � )    � .    � 7    � 8    � 9    � :    � <    � =    � ?    � @    � B    � C    � E    � H    � M    � V    � W    � X    � Y    � \    � ]    � `    � b    � e    � f    � g    � h    � i    � j    � k    � l    � l     n    o    p    s    x    �    �    �    �   	 �   
 �    �   S�e��a�1J   �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �     �   ! �   " �   # �   $ �   % �   & �   ' �   ( �   ) �   * �   + �   , �   -    . 	   / 
   0    1    2 )   3 *   4 +   5 ,   6 ,   7 -   8 .   9 /   : 0   ; 0   < 1   = 2   > 3   ? 5   @ 9   A     B  �   C  �   D  �   E  �   F  �   G  �   H  �   I  �   J  �   K  �   O��>-�e��E�  L  �   M  �   N  �   O  �   P :   Qnnnn���@�����@@@@@@@      X      ��������������  ���� �P    �  �      @������  ����                                                                                                                                                                                                                                                                                                                                                                                          !%=�N;�x�7                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   �    � [�D         !N7�  D               �  `                                                                                                                                                                                                                                                                                                                                                                                                                                                                         	�y�����8Y H                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  
�s�Xo   �@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   �`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   �                            0     p      0�����@����@�����\���������@@@@@@��������@@�����@@@@@            �������������   ��������        \���         �@                \���     �` �0                                                                                                                  p           7������@@@@\����@@@@@          7����@@@@@@\����@@@@@          7��������@@\����@@@@@                                                                                                            �ʊ��0��9G#�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �s�Xo   �@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   �`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   �  �����������@@@@@@@@@@@@@@@@@@@@@@@  �                              �      @ @           (                                                   �a�@������@����������@@@            ����  �s�TU�   �                                                  �>n�  С0�Y �                                                                                                                                                                                                                                                  }���������                                                                                                                                      �>n�                                                                                                                                                                                                                                                                                                                                                                                     �s�XO =Y�P                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �s�Xo   �`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo   �    �� �>n�          �>n�  � �������@@@@@@@@@@@@@@@@@@@@@@@         @�s�ݾ�  .�M��           
~6O   �>n�         �s����                          �   �                                �                                       �                ��������@@\����@@@@@  \@@@@@@@@@@@@@@@@@@@ ����^�������@@@\����@@@@@                             :@        y �-^�� �  �      
        	    ����@@@@@@  �   	.� ��`          	�    ���@@@@@@@  � z   �zz   	��K   l    !��|��t_�       @ 	�    ������@@@@ K �    ������  ��   	���   d  F       @ 
    �������@@@ � �    ���   
&��   d         @ 
E    �������@@@ � �    ���   
c�.   P          
{    ��������@@ . � # �����(:EUh�   
��w   P         
 
�    ��������@@ w �  ������   
���   l           
�    ���������@ � �    �������  ��   
� m�3   l               ���������� 	3   "jz o��� `k��    �������   ��   ' m�{   H           M    ���������@ 
{ !  	   d m��   H           u    ���������@ � !  	   � m�   l           �    ����@@@@@@      ��  �   � m�_   H           �    ���������� _ !  �!   � m��   H           �    ���������@ � !  �!    m�     P  
        $    ������@@@@    # 	 #.   < m�  �   
          #���wT��-� 	?     �   	L��=  �   
         	]       	n��    �           	      ��   	���    @ @�  \ @ ������ ������ \����    \����      	��� \������ \���� \��� Ö����� Ö�����`�� Ö�����`ւ����� Ö�����`��ւ����� ㉔��`ٖ��� 
㉔��`�� ㉔��`ɣ���� ㉔��`��ɣ���� 	ȅ������� ȅ�������`�� ȅ�������`ւ����� ȅ�������`��ւ����� ⨔��� 遗�ĉ������ \���� \���������� \����������� \������������ \������������ \������ \�� Y_ \�� �/ \������ a/   $Ge�ʠ�֪�� y/ �� __ � � \��� � ��  	\�������� 
\��������� �\����@@@@@@@@@@@@@@@\����@@@@@m������      \@@@@@@@@@@@@@@@@@@@         %\����@@@@@@@@@@@@@@@   �                                                               \����@@@\����@@@\����@@@@@@@@@@@@@@@\����@@@@@\����@@@@@@@@@@@@@@@\����\����@@@                                                                                                                                                                                             @@@@@@@   Ö�����@���  %��^d�D�--�@◖��Ɖ��@����@��� 
@@@@@@@   ◖������@���� @@@@@@@   Ձ�� 
@@@@@@@@@   @@@@@@@   Ձ�� 
@@@@@@@@@ 䢅� @@@@@@@   Ձ�� @@@@@@@@@ դ���� @@@@@@@   ������`������ @@@@@@@@@ і�@����  @@@@@@@   \ @@@@@@@@@ ◖������@������ @@@@@@@   �`������k@\����k@\���� F@@@@@@@@@ 
���@������ 	@@@@@@@   ׁ��@����k@\������ @@@@@@@@@ ���@��������@���� @@@@@@@   Ձ��k@\���� @@@@@@@@@ ��Ɩ��  @@@@@@@   
Ö�����@KK @@@@@@@@@ ׁ������  @@@@@@@   	\����@KKK @@@@@@@@@ 
ׁ��@扄�� @@@@@@@   �`����k@\�  &�a��QU����k@\��k@\������ @@@@@@@@@ ׁ��@ȅ���� @@@@@@@   �`����k@\��k@\��k@\������ @@@@@@@@@ 
ז���@≩� @@@@@@@   �`�� @@@@@@@@@ 兙�����@◁�� @@@@@@@   �`�� @@@@@@@@@ ׁ��@ȅ���� @@@@@@@   �`���k@\��� @@@@@@@@@ Ӆ��@ԁ���� @@@@@@@   �`��� @@@@@@@@@ 
㖗@ԁ���� @@@@@@@   �`��� 
@@@@@@@@@ ֙���������  @@@@@@@   \��������k@\���������\����@@@@@@@@@@@@@@@                                                                                                                                                '�S��p_rU�/�7                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  (�s�Xo   �  ������������K�@@@@@@@@@@@@@@@@@@@@�                                  �   '   @ @   0                                                            �a�@������@����������@@@            ����  �s�TU�   �    (                                               ���  �j�� �                                                                                                                                                                                                                                                  )��&�an�ecr�                                                                                                                                  @   @ ���                                                                                                                                                                                                                                                                                                                                                                                     *�s�X� -�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   +�s�Xo   �`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ,�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   -�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   .�s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   /�s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   0�s�Xo   �     �� ���         ���  � ���������K�@@@@@@@@@@@@@@@@@@@@�   0     ��s�V�� "�Ф�                   ���         �s�]2�                           �   �                                �                                      �                                                                                                                                                                                                                                                                                1g^E�HF����E�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  2�s�Xo   �@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   3�s�Xo   �`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   4�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   5�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   6�s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   7�s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   8�s�Xo   �  C�������@@@@@@@@@@@@@@@@@@@@@@@�s�dG         @@�������  \������@@@    �   \������@@@                      ��������@@@@@@@@@@@@@@@@@@@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@    �     	P  `                 @@@@@@@@@@@@@@@@@@@@                                 ������@@@@@@@@@@@@@@@@@@@@@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@    �   7  `  @                 @@@@@@@@@@@@@@@@@@@@                                                                                                                                     9N�Ǉ��@�ghrL                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  :�s�Xo   �@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ;�s�Xo   �`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   <�s�Xo   �                                                                                                                                                                                                                                                                                                                                                      �          @      �� @                              @@��         �        \�������@@      5         <   @   �������������  @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  =f>�j*�3]� @@@@@@@@@@@@@@             ������@@@@��������@@�������@@@��       �  '�                      @�����   %            .K��"         .K��"                                           �   �                 �            `              �                                                                                                                                                                                                                                                                                  >�Z.}Rn�O|G�                                                                                                                                                                                                                                                                                        K��                      ���������@�                                                 @@@@@@@@@@@@@@@@@@@@@�����������                                                        (�fɫ                % %        ��  � ����������@��  ?�C�ȗ&&�P�^������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �����@@@@@@����@@@@@@                               2 �          �         % % %                                                           ��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ �����@@@@@@����@@@@@@    �                         2 �          �         % % %                                                          ��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                                                       @�E�P�sj�#�                                                                                                   ���������@@     p   !   �   !               @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �������������        .K��"                                  @@@@@@@@@@                                                     ��������@@��������@@@@@@@@@@@@�       �@@@@@@@@@@@@@@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@��������������������������������������@@@@��������@@�������@@@@@@@@@@@@@@@@@@                                  Asamre�E�}���@@                 �������@@@��������               ��@@@@@@@@�                                              @      �� @                              @@�h         �        \�������@@        5         <   @   �������������  @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                                           ��       �  '��                     @�����   %            	�Fdl         (�ہ                                           �   �                 p            `                 Bj��w�=��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  C�s�Xo   �`                                         /S���                      ������@@@@�                                                 @@@@@@@@@@@@@@@@@@@@@�����������                                                        ŧ��                % %        0��  � p������@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �������@@@@������@@@@                                                                                                                      �������@@@@������@@@@       D�#�+ʷ��^�                                                                                                               �������@@@@������@@@@    d                                                 %                                                                                                                                                                                                                  ���������@@     p   !   �   !               @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �������������  E�@����fo�        	�Fdl                                 ��@@@@@@@@          �������������                 ��������@@@     p   !   �   !               @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �������������        ۈ$y                                 �����@@@@@  d      �������������                 ��������@@@     p   !   �   !               @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �������������        J���                     S            ���@@@@@@@          �������������                F�}Y���*IA~]   ���������@@     p   !   �   !               @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �������������        !&�H                     �            ����@@@@@@          �������������                 ���������@@     p   !   �   !               @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �������������        &՞�                                 �����@@@@@  d      �������������                 ���������@@     p   !   �   !               @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  G�ʲ�Y��l�@  �������������        (�ہ                    5            �����@@@@@  d      �������������                              ������@@@@��������@@@@@@@@@@@@�������@@@@�������@@@@@@@@@@@@@�������@@@@�������@@@@@@@@@@@@@�������@@@@��������@@@@@@@@@@@@�������@@@@��������@@@@@@@@@@@@�������@@@@��������@@@@@@@@@@@@�       �@@@@@@@@@@@@@@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@�������������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                                @@                 �������@@@��  HI�lo��=�[�6������               ��@@@@@@@@�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                I�s�����rh�@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  J�s�Xo   �@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   K�s�Xo   �`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   L�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   M�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   N�s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   O�s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   P�s�Xo   �  ������������@@��������@@@@@@@@@@@@�   p                                    ]@ @                                               `                �a�@������@����������@@@            ����  �s�TU�   �                                                      �   �WM�D �                �WM�D �                        �WM�D                                                                                                                                                                                            Q[��xu���X�8                                                                                                                                      0@�         ���                                                                 �                                                                                                                                                                                                                                                                                           R�s;�R���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  S�s�Xo   �`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   T�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   U�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   V�s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   W�s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   X�s�Xo   �     �� 0@�              �   � ���������@@��������@@@@@@@@@@@@          @]�s��/C  .�M��                   0@�          �s��/u                           �   �                                �                      .K��"            �                \            0@� `0@� 0                                           '      '      �        @  �                  �0@�          @�������       �                                                                0@� P                          YDl�_�� S0m                                                                             G�0@� @                                      �               �                                                        ���     ]                                                                                                                                                                                                                                              ��                                                            Z�rޓ~��,�                                                              �                           �@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@        ��� �      �                                                                                                                                                                                                   [���V�W1�T                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  \�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ]�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ^�s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   _�s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   `�s�Xo   �    �  0@�             �   �@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                                                                                                                                                                                                                                                                                          a�ނ��ϳt�H                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  b�s�Xo   �@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   c�s�Xo   �`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   d�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   e�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   f�s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   g�s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   h�s�Xo   �  ����������@@@@��������@@@@@@@@@@@@�                                0      ]@ @                                               �                �a�@������@����������@@@            ����  �s�TU�   �                                                      �   �A�n �                �A�n �                        �A�n                                                                                                                                                                                            i�(;����Ro                                                                                                                                       :�|��         "la�!                                                                                             d                                                                                                                                                                                                                                                           j�{)3�KS&ˠ                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  k�s�Xo   �`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   l�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   m�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   n�s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   o�s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   p�s�Xo   �     �� :�|��              �   � �������@@@@��������@@@@@@@@@@@@          @]�s���� .�M��                   :�|��          �s��ư�                           �   �                                �    �t              	�Fdl            �                j�           :�|�� �:�|��                                     "      '      '      �        @  �                  q:�|��          @�������      �                                                                :�|��           @                qC�1^��rb-                                                                            C�:�|��                                       p               q                                                        ���     ]                                                                                                                                                                                                                                             �M>�0                                                            r�r��e`L-!6-                                                                                          d                           �������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@               "la�! �      �                                                                                                                                                                                                                                                   s�W�ʸ��vƛ                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   t�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   u�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   v�s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   w�s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   x�s�Xo   �    �  :�|��             q   �������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@@@@@@@@@�@���������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������M}����}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@@@@@@@@  y7y,!���%(�+@@@����@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������M}����}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                                                                                                                                                                                                                                                                                                                            z�ڔ�Y&m���:(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  {�s�Xo   �`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   |�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   }�s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ~�s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   �  ����������@@@@�������@@@@@@@@@@@@@�                                0      ]@ @                                               �                �a�@������@����������@@@            ����  �s�TU�   �                                                      �   Ұ�
� �                Ұ�
� �                        Ұ�
�                                                                                                                                                                                            �L�kx#��	Ҙ                                                                                                                                      (1٭�         ���                                                                                             d                                                                                                                                                                                                                                                           ��{0i`���0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��s�Xo   �`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   �     �� (1٭�              �   � �������@@@@�������@@@@@@@@@@@@@          @]�s���E� .�M��                   (1٭�          �s���                            �   �                                �    �t              ۈ$y            �                m�           (1٭� �(1٭�                                     "      '      '      �        @  �                  q(1٭�          @�������      �                                                                (1٭�           @                �B1\�oO��eR��                                                                            C�(1٭�                                       p               q                                                        ���     ]                                                                                                                                                                                                                                             ���                                                            ��r�������3�                                                                                          d                           �������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@               ��� �      �                                                                                                                                                                                                                                                   ��W�ʸ��cӷ]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   �    �  (1٭�             q   �������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@������@@@@@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@ؤ�@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�������@@@@@@@@@@@@@@@@@�@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@¨���@�  ��O�������$�������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�������@@@@@@@@@@@@@@@@@�@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@¨���@���������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�����@@@@@@@@@@@@@@@@@@@�@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@ŧ�������@Ʉ@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ���{>2�$�[n�@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@��������@@@@@@@@@@@@@@@��@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@偙����@������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@���������@@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@ؤ�@��������@@  ���T��[��
D5@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@������@@@@@@@@@@@@@@@@@@�@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@҅�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���������@@@@@@@@@@@@@@@�@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@¨���@י������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �:�qL�S;�Sav@@@@@@@@@@@@@@@@@@�������������@@@@@�@���������@@@@@@@@@@@@@@@�@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@¨���@���������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�������@@@@@@@@@@@@@@@@��@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@ŧ�������@Ʉ@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@����������@@@@@@@@@@@@  ��V���F��ȯ�@��@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@م������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@����������@@@@@@@@@@@@��@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@��������@@@@@@@@@@@@@@@��@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��h�H}?N���;@@@@@@@@@@@�������������@@@@@@\@ֆ����@ŧ�@ā��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@��������@@@@@@@@@@@@@@@��@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                                                                                                                                                                                                                                                                                     ��4K�z��*���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��s�Xo   �  ����������@@@@�������@@@@@@@@@@@@@�                                0   '   ]@ @                                               �                �a�@������@����������@@@            ����  �s�TU�   �    (   	                                                �   ʬn� �                ʬn� �                        ʬn�                                                                                                                                                                                            ���:��TA8                                                                                                                                      .�;     0   0 3���                                                                                             d                                                                                                                                                                                                                                                           ��{"k�F}pp                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��s�Xo   �`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   �     �� .�;              �   � �������@@@@�������@@@@@@@@@@@@@           @]�s��1	� .�M��                   .�;          �s��J��                           �   �                                �    �t              J���            �                �           .�; �.�;               S       S               k      '      '      �        @  �                  q.�;          @�������      �                                                                .�;          @                �C�0)�(�:�=                                                                            C�.�;                                       p               q                                                        ���     ]                                                                                             S                                                                                                                                                ��0                                                            ��r��D��H�	                                                                                          d                           �������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@               3��� /�      �                                                                                                                                                                                                                                                   ��W�ʨ�	`�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ��s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   �    �  .�;             q   �������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\@@�������z@�������@�@�����@���@����@���@��������@@@@@@@@@@@@@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@  ��"L�M�G#Ɣ��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@���@������M}Ö�����@���@◖��Ɖ��@����@���}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@����@����@@@@@@@����M\����]@���M��]@���M�]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M}◖������@����}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��jN�F���@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@����@���@@@@@@@@����M���]@���M\]@������MM\]]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M}і�@����}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@����@������@@@@@����  �z��{����pM\���]@���M�]@���M\����]@�����M�@������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������MM\����@�]@M\����@`�]]@����M\���]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M}◖������@������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@����@�������@@@@����M\�����]@���M��]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��6Ǉ%���S��@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@���M\������]@������MM\������]]@���M�]@����M\���]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M}���@������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@����@�������@@@@����M\�����]@���M��]@���M\����]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������MM\��  ��� �i(�S{�d��]]@���M�]@����M\���]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M}���@��������@����}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@����@��������@@@����M\����]@���M��]@����M\���]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@���M\���]@������M\���@}Ö�����}@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �ڑ=|&tթ�u@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@}Ö�����`��}@}Ö�����`ւ�����}@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@}Ö�����`��ւ�����}@}㉔��`ٖ���}@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@}㉔��`��}@}㉔��`ɣ����}@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@}㉔��`��ɣ����}@}ȅ�������}@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@}ȅ�������`��}@}  ���,��N
�g�2�ȅ�������`ւ�����}@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@}ȅ�������`��ւ�����}@}⨔���}@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@}遗�ĉ������}]@������M}Ö�����@KK}]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M}��Ɩ��}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��]����3�A�@@@@�������������@@����@��������@@@����M\����]@���M��]@����M\���]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@���M\����]@������M\����@\����������@\�����������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@\������������@\������������@\������]@������M}\����@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@KKK}]@������M}ׁ������}]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �L��K}w$z]�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@����@���������@@����M\���]@���M�]@���M\��]@�����M�@����]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������MM\��@���]@M\��@���]@M\������@���]]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M}ׁ��@扄��}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���  �P�D��m~=�9�����������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@����@����������@����M\���]@���M�]@���M\��]@�����M�@����]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������MM\��@���]@M\��@����]@M\������@���]]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M}ׁ��@ȅ����}]@@@@@@@@@@@  ��leF �Na�p}@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@����@���������@@����M\���]@���M�]@���M��]@�����M�@��]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M}ז���@≩�}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����������  �)h�K�I�g {����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@����@���������@@����M\���]@���M�]@���M�]@�����M�@��]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M}兙�����@◁��}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ����@�~] 2@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@����@����@@@@@@@����M\���]@���M�]@���M\���]@�����M�@���]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������MM\���@`�]]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M}ׁ��@ȅ����}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@  ���$�N�Ԏ'O�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@����@����������@����M\���]@���M�]@���M��]@�����M�@���]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M}Ӆ��@ԁ����}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �0�����pb�֦@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@����@���������@@����M\���]@���M�]@���M��]@�����M�@���]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M}㖗@ԁ����}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@����@����  ���Z��z#�O���@@@@@����M\����]@���M��]@����M\���]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@���M\��������]@������M\��������@\���������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@������M}֙���������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �88edf^�#@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����������������z@����@����M\����]@���M\]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@����@����M\����]@���M��]@������M}䢅�}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@����@����M\����]@���M�]@�����M������@������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@������M}դ����}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@  �<6�_�q�"h#b�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��������������������z@������@���M��������]@����MM\��@\������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                                                                                                                                                                                                              �m���!R�η�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   �  ����������@@@@��������@@@@@@@@@@@@�                                0   ?   ]@ @                                               �                �a�@������@����������@@@            ����  �s�TU�   �    @   
   8                                            �   �/$�Z �                �/$�Z �                        �/$�Z                                                                                                                                                                                            ���^KZ8��_�\                                                                                                                                      �]-�     `   ` 9�A��                                                                                             d                                                                                                                                                                                                                                                           {.$��0��`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  És�Xo   �`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ĉs�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ŉs�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   Ɖs�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ǉs�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ȉs�Xo   �     �� �]-�              �   � �������@@@@��������@@@@@@@@@@@@         8 @]�s��w
� .�M��                   �]-�          �s����                           �   �                                �    �t              !&�H            �                @           �]-� ��]-�               �       �               �      '      '      �        @  �                  q�]-�          @�������      �                                                                �]-�          @                �B4����s�g�=                                                                            C��]-�                                       p               q                                                        ���     ]                                                                                             �                                                                                                                                                ��0��                                                            ʉr��4�p�T��                                                                                          d                           �������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@               9�A�� _�      �                                                                                                                                                                                                                                                   ˙W��P�&W?w                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ̉s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ͉s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   Ήs�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ωs�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   Љs�Xo   �    0�  �]-�             q   �������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@����MP����@P���@P������@P�������@P�������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@P��������@P��������@P���������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@P����������@P���������@P���������@P����@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@  �E�b���f-4�C�@@@@@@@@@@@P����������@P���������@P������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���������@@����M}ǉ������@Ö���������@����@`@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@����������|�����K��}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP����]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP���]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@  �R:I�� �|�>C�@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\���]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP�������]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP�������]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP��������]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@  ��h��?�h%֥@@���MP��������]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP���������]@����M\���]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP����������]@����M\���]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP���������]@����M\���]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP���������]@����M\���]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@  ��E�h�gX3��@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP����]@����M\���]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP����������]@����M\���]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP���������]@����M\���]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP  գ /Ȱ���3N�������]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP����]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP�������]@����M\����]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP�������]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��e�c���Tn%@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP�������  כ��I���N���]@����M\����]@���M����]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@���M���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP����]@����M\����]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP�]@����M\���]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP�������]@����M\����]@���M���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �X�t����\�-@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP���]@����M\����]@���M���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP����]@����M\����]@���M�]@�����M�}��}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@���M���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP�������]@����M  �f�N����7~�\����]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP����]@����M\����]@���M���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP�����]@����M\����]@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@@@@@@@@���MP������]@����M\����]@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���  ڞi�QR�2�k�z����������@@@@@@@@@@@@@���@@@@@@@@���MP�������]@����M\���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@�����M�������]@����M����@������M�����]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\@ǅ�@���@����������@��@���@�������@����@@@@@@@@@@@@@@@@@@@@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\````````````````````````````````````````````````  ��Eo����&�x````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���MP����]@�����M}�}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@��@@@@@@@@@����MP���@~@}\}]@����M�������@���MP�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@����MP����]@���MP������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@����@@@@@@@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����������  ܵW�L�f:�썢����@@@@@@@@@@@@@������@@@@@���MP�������]@�����Ml���MP���@�@��]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���MP����]@�����Ml���MP���@��@��]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���MP������]@�����Ml���MP���@��@�]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���MP�������]@�����MP������]@@@@@  �:��Ck�è>�1@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���Ml���MP������]]@�����MP�������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���Ml���MP������]]@�����M����]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���MP������]@�����M�}����������������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@����@@@@@@@���M��������]@����MP��������@P������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@  ޢ��.�����7w@@@@@@@@@@@@@@@@@@@@@@}��������}@P���@}@}@}@}@P����@P������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@P������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���MP�����]@�����Ml���MP������@�@�]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@��@@@@@@@@@����MP�����@\��@}@}]@����M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���MP������]@�����Ml���MP������@��@��]]@  ߈��V��$�rT@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���������@@�����MP�����]@����M�������]@������MP������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@�������M\������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\@È���@��  ��c�%���B㢅@������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���MP�������]@�����Ml���MP��������@���@��]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@��@@@@@@@@@����MP�������@\��@}\���}]@����M���������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@�����M�������]@����M�������]@N@@@@@@@@@@@@@@@  �<�y�kq����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@������M}◖��@��@���@\���}]@�������M\������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\@È���@��@���@���������@��@����������@��@���@�����@@@@@@@@@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@��@@@  �_���Ϫ�bK�@@@@@@����MP������@~@`�]@����M������@���MP�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@�����M\����]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@����@@@@@@@���M��@����MP������@~@�]@����M������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@���MP�������]@�����M\����]]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@��������@@@����MP����]@���MP������aP����aP�������]@N@@@@@@@@@@@@@  ����+vV/d@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@������MP�������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\@È���@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\@ׁ��@�������@\a@@@@@@@  �M��g�Y���m@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@��@@@@@@@@@����MP�������@~@}@}]@����M���������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@�����M�������]@����M�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@������M}ׁ�������@�������@�������}]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@�������M\������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��5 
�0$ڏ_�@@@@@@@@@@@@@@@�������������a\@ą�����@����@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@��@@@@@@@@@����MP�������@~@}\������}]@����M����@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@���M��������]@����MP�������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\@È���@ׁ��@���������@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���MP���  ����D��de���]@�����M}�}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���MP�]@�����M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���������������������z@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���MP�]@�����MP�@`@�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@��@@@@@@@@@����Ml���MP�������@P�@�]@~@}a}]@����M����@N@@@@@@@@@@@@@@@@@@@@@@@@@  �`�e���xlW4@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@������M���������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@��@@@@@@@@@����Ml���MP�������@P�@�]@~@}@}]@����M����@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@������M��������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���MP�������]@�����MP�������@\����@}a}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����������������������z@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ���]�v\�+�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���MP�������]@�����MP�������@\����@P����]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@�������@@@@���M}����}]@����MMP�������]@MP������]]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@������Ml���MP������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@��@@@@@@@@@����Ml���MP������]@\��@�]@����M���������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �wuh���ߐ�錥@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@�����M�������]@����M�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@������M}晖��@ׁ��}]@�������M\������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\@È���@���@Ձ��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\````````````````````````````````````````````  ��ji��rİ�2�````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\@�������@�������@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@��@@@@@@@@@����MP�������@~@}@}]@����M���������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@�����M�������]@����M�������]@������M}���@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@����@�������}]@�������M\������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������  �=B�w�u���w�������a\@ą�����@�������@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@��@@@@@@@@@����MP�������@~@}\����}]@����M������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@���MP�������]@�����MP����]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\@Ö��@���@◖��@����@�@��@@@@@@@@@@@@@@@@@@@@@@@@@@  �=C\M���SU%)@@@@@@@@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\@ǅ�@���@�����@����@����@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���MP������]@�����Ml���MP��������@���@�]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���MP������]@�����Ml���MP��������@���@�]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������  홾�wI�I��˙�a\@���@�@������@���@����@�����@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���MP����]@�����M}�}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���������@@������M�����]@������MP�������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���MP������]@�����M}�}@\���@P�������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@����M����a��������]@���MP������]@@@@  �9OrC�]��T\�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@�����M�������]@����M������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@����M����a��������]@���MP������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@�����M�������]@����M���������@�����M�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@����M�������]@������M}���@����@���@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@  ��x�b��0ח�@@@@@@@@@@@@@@@@@@@�����}]@�������M\������]]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\@Ö��@���@���������@����@���@������@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���MP����]@�����M}�}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@�������@@@@����MP����]@������M����a��������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@���MP������aP����aP�������]@N@@@@@@@@@@@@  �Tg3a�p�Q@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@������MP�������]@�����MP������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@������M\���]@�������M\����]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\@Ù����@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\````````````  �fT��������````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���MP���]@�����MP�������@\����@P�������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@\����@}K���}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@����@@@@@@@���M��������]@����MP����@P������@P������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@P������@P���@P��������@P��������@N@@@@@@@@@@@@@@  �	������ҥ�@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@P���������@P����������@P���������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@P���������@P����@P����������@P���������@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@P������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\@ㅙ������@@@@@@@@@  �5�az��Xw�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\````````````````````````````````````````````````````````````````\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\@م����@���@���������@����@��@���@�����@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@����@@@@@@@����M����a��������]@���MP������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@����M\����]@�����M\���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �j\��2�2���@@@@@@@@@@@@@@@@@@@�������������a\@⅕�@�@����������@�������@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���������@@�����M�������]@����M�������]@������M}◖��@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@����}@\����@P����@\����@}���������@����}@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@\����@P�������@\����@P�������@\����@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@}K  �	zX�Td�مW���}]@�������M\����]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\@ř����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������a\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\a@@@@@@@@@@@@@@@@@@  �"�;�|�Q�@@@@@@@@@@@@������������������z@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@��@@@@@@@@@����MP�������]@����M���������@�����M�������]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@����M�������]@�������M\������]]@a\@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@��������@�����@@@@@@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@���MP������  ��.C�Xü˂���]@�����M}�}]@a\@���@������@��@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@�����@@@@@@\a@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@����@@@@@@@���M��������]@����M}@@@@}@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@�}������������������������������}@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@�}�����������������������������������������N@@@@@@@@@@@@@@@@@@@@@@@@@  �t��h�<J|���@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@�������������������������������������������N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@������������}@�}��������}@��������@\@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@�}��������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                                                         �c!��6�D"���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��s�Xo   �@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   �`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��s�Xo   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo     ����������@@@@��������@@@@@@@@@@@@�                                0      ]@ @                                               �                �a�@������@����������@@@            ����  �s�TU�   �                                                      �   ��%�� �                ��%�� �                        ��%��                                                                                                                                                                                            ��U��Gs@���                                                                                                                                      ��I)         ?G�t                                                                                             d                                                                                                                                                                                                                                                           �{'�^I�j�P                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �s�Xo   `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo       �� ��I)              �   � �������@@@@��������@@@@@@@@@@@@          @]�s���� .�M��                   ��I)          �s���                            �   �                                �    �t              &՞�            �                ;`           ��I) ���I)                                     "      '      '      �        @  �                  q��I)          @�������      �                                                                ��I)           @                	B�ǂ���dK{=                                                                            C���I)                                       p               q                                                        ���     ]                                                                                                                                                                                                                                             ��}Ր                                                            
�r���"M��:�                                                                                          d                           �������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@               ?G�t �      �                                                                                                                                                                                                                                                   �W�ʸ���b�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo      �  ��I)             q   �������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@Ć�������M\��]@������M\���]@������M}�����}]@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���������@@M}ǉ������@Ö���������@����@`@����������|�����K��}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa```````````````````````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@ׁ����  S�Iu�Yt�=�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa```````````````````````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ŕ���ׁ���@@@@@@@��@@@@@@@@@@@@@@@@@@������M}��������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@ׁ��@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ŕ���ׁ���@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �H"�� k�U�̀@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@ׁ��@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@���@����@����@��@�������@�������@���������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@ć�����@@@@@@@@@@@��@@@@@@@@@@@@@@\@@@�������M}������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���ĉ�@@@@@@@@@@@@@@@@@@@@@@@@@@\@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���≩�@@@@@@@@  F�d[t�u��$�@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���ĉ�@@@@@@@@@@�@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@aa@���������@���@�������@���������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@��@M������Ml����Mä����]z@l����M������]]@~@\����]^@@@@@@@@@@@@@@@@@@@@@@@@@  ����#�f	G�f@@@@@@@@@@@@@@@@@@�������������@@@@@@@ׁ��@~@}@}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@ׁ��@~@l���Ml����Mä����]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@\����@~@\��^@@@@@@@@@@  `,'b�y��r	@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                                                                                                                                                                                                                                                                                                                                           �P�MU[ϲp                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �s�Xo  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo    ����������@@@@��������@@@@@@@@@@@@�                                0   �   ]@ @                                               �                �a�@������@����������@@@            ����  �s�TU�   �    �      �                                            �   Ҧ��X �                Ҧ��X �                        Ҧ��X                                                                                                                                                                                            L.T����i7[                                                                                                                                      26�    p  p ,�	6                                                                                             d                                                                                                                                                                                                                                                           �z�.��'��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �s�Xo  `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �s�Xo  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �s�Xo       �� 26�              �   � �������@@@@��������@@@@@@@@@@@@         � @]�s���O  .�M��                   26�          �s��x�                           �   �                                �    �t              (�ہ            �                Z            26� �26�              5      5              @      '      '      �        @  �                  q26�          @�������      �                                                                26�          @                !C$1�x���                                                                            C�26�                                       p               q                                                        ���     ]                                                                                            5                                                                                                                                                ���@                                                            "�r��d��v3�                                                                                          d                           �������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@               ,�	6o�      �                                                                                                                                                                                                                                                   #�W����?,S�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   $�s�Xo  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   %�s�Xo  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   &�s�Xo  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   '�s�Xo  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   (�s�Xo      ��  26�             q   �������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@Ć�������M\��]@������M}�����}]@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���������@@M}ǉ������@Ö���������@����@`@����������|�����K��}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa```````  )3C��&�C��````````````````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@◖��@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa```````````````````````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@���������@@��@@@�@@@@@@@@@@@@@����@@@@������M�������]@������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  *�;��	���r`@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa```````````````````````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@Ô�@ׁ��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa```````````````````````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ŕ���ׁ���@@@@@@@��@@@@@@@@@@@@@@@@@@������M}��������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�����@@@@@@@@@@  +�&��)�m�)$�@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�������@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�������@@@@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�������@@@@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@������@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ,:ܢ��vX�+Cb�@@@@@@@@@@@@@@@@@@�������������@@@@@�@���������@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���������@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@����������@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�����������@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@����������@@@@@@@@@@@@  -(?E�d�:�t@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@����������@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�����������@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@����������@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  .߹�0I]�����@@@@@@@@@@@�������������@@@@@�@�������@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ŕ���ׁ���@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�������@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�������@@@@@@@@@@@@@@@@@@@@@@  /����7�c6��?X@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�������@@@@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@������@@@@@@@@@@@@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���������@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���������@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  0��hV�`mP�@@@@�������������@@@@@�@����������@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�����������@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@����������@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@����������@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@��@�@  1JՐ�W���mA�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�����������@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@����������@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�������@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���  2����ܯ+j�f����������@@@@@������@@@@@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@ؤ�@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�������@@@@@@@@@@@@@@@@@�@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@¨���@י������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�������@@@@@@@@@@@@@@@@@�@@@@@@��@�@@@@@@@@  3��FC�P�I���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@¨���@���������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�����@@@@@@@@@@@@@@@@@@@�@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@ŧ�������@Ʉ@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@��������@@@@@@@@@@@@@@@��@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����������  4H��Bh(�#�����@@@@@@\@偙����@������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@���������@@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@ؤ�@��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@������@@@@@@@@@@@@@@@@@@�@@@@@@��@�@@@@@@@@@@@@@@@  5�]�h�*J4���y@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@҅�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���������@@@@@@@@@@@@@@@�@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@¨���@י������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���������@@@@@@@@@@@@@@@�@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@  6?Cb�S<�nNk��@@\@¨���@���������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�������@@@@@@@@@@@@@@@@��@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@ŧ�������@Ʉ@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@����������@@@@@@@@@@@@@��@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@م������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  7�j�dpn��SB��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@����������@@@@@@@@@@@@��@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@��������@@@@@@@@@@@@@@@��@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@\@ֆ����@ŧ�@ā��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@����  8�γ����R�����@@@@@@@@@@@@@@@��@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@��������@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@⣙���@����@��ɢ@``````````````````````````````````````````````````K@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@Ĥ�����@@@@@@@@@@@��@@@@@@@@@@@@@��@�@�������M}������}]@@@@@@@@@@@  9SB����v{��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@Ė���@@@@@@@@@@@@@��@@@@@@@@@@@@���@�@�������M}����}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@@@@@@@@@@@  :󸅫������ǘ@@@@@@@@@@@@@@@@@@@���@�@�����@�������M\������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@�������M\������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�m�����@@@@@@@@@�@@@@@@@@@@@@@���@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�m������@@@@@@@@�@@@@@@@@@@@@@���@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�m�����@@@@@@@@@�@@@@@@@@@@@@@���@�@���M��]@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ;�4�֒�x7�	�S@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�m��������@@@@@@�@@@@@@@@@@@@@���@�@���M�������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�m�����@@@@@@@@@�@@@@@@@@@@@@@���@�@���M���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�m�����@@@@@@@@@�@@@@@@@@@@@@@���@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@Ħ����@@@@@@@@@@@@��@@@@@@@@@@@@���@�@�������M}�����}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@@@@@@@@@@@@@@@@@@  <��Z��;�Z�@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@ă����@@@@@@@@@@@@��@@@@@@@@@@@@���@�@�������M}�����}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  =:�0�+��u@@@@@@@@@@@@@@@�������������@@@@@@aa@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@Ć�@@@@@@@@@@@@@@@�@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@Ӗ���@����������@``````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�Ⅳ��ׁ��@@@@@@@@��@@@@@@@  >��!d����Ԟ2@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�Ù���Ƣ���@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@������@@@@@@@@@@@@@@@@@@@@@@@����@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉��ȅ����@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ?�j(.��\�r�@@@@@@@@�������������@@@@@�@㉣��@@@@@@@@@@@@@@@@@@@@@@@@����@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉��ׁ���@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉��ׁ���㙅�@@@��@@@@@@@@@@@@@@  @��!)��ϻ#t�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉���م�@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉��㙁����@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  Aa�k��܈����@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�⣁��ׁ��@@@@@@@@��@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ŕ�ׁ��@@@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@⣙���⣁��@@@@@@@@@@@@@@@@@@@���@�@@@@  B�ev:�]oL���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉��ā��@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@¤����@@@@@@@@@@@@@@@@@@@@@@�����@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@Ӆ�@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������  Cdf��26��� ��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�Ó�����Ƣ���@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ɕ�ん�����@@@@@@��@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  D[@b�K&���`�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ǅ�ř�ɕ��@@@@@@@��@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�╄ׇ�Ԣ�@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@����@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������  E�-M�o�_ؓ��@@@@@�@��������@@@@@@@@@@@@@@@@@@@@@@���@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���Ʉ@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���@@@@@@@@@@@@@@@@@@@@@@@@@@����@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  F�5yH��=�ZR�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@Ö��������@�����@``````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ん�����@@@@@@@@@�@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@ԉ��@���������@````````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@��  G�]�K��sَ�w�@@@@@@@@@@@@@@@�@@@@@@@@@@@@@@@@@@@�}��}@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@���@偙������@`````````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ׁ��Ֆ@@@@@@@@@@@�@@@@@@@@@@@@@@��@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ׁ��ւ����@@@@@@@�@@@@@@@@@@@@@@��@�@���M���]@@@@@@@@@@@@@@@@  Hʭ!��j����qy@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@ħւ����@@@@@@@@@@�@@@@@@@@@@@@@@��@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@ħֆ����@@@@@@@@@@�@@@@@@@@@@@@@���@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@ħم�@@@@@@@@@@@@@�@@@@@@@@@@@@@���@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�Ӗ�������@@@@@@@@�@@@@@@@@@@@@@���@�@���M����]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@  I�b8���̺p0�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ז���≩�@@@@@@@@�@@@@@@@@@@@@@@��@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�兙�◁��@@@@@@@@�@@@@@@@@@@@@@@��@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�Ö��@@@@@@@@@@@@@�@@@@@@@@@@@@@@��@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�Ӆ��ԁ����@@@@@@@�@@@@@@@@@@@@@@��@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@  J+f n(o�dNP�@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�㖗ԁ����@@@@@@@@�@@@@@@@@@@@@@@��@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ׁ��扄��@@@@@@@@�@@@@@@@@@@@@@@��@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ׁ��ȅ����@@@@@@@�@@@@@@@@@@@@@@��@�@���M�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@  K�3lJ����}��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ą�����Ɩ��@@@@@@�@@@@@@@@@@@@@@@@@@@}Ö�����}@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�Ɩ��@@@@@@@@@@@@@�@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  L</�-�n�7�ʈ@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@י�����@������@````````````````````````````````````````````````````@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ׇ�⣢@@@@@@@@@@���@@@@@@@@@@@@@@@@@@Ֆ֗�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@і�Ղ�@@@@@@@@@@@@@@@@@@@@@@@@@��@@@֥�����Mׇ�⣢z���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa\\\\\\\\\\\\\\\\\\\\  M��m�2i��^O�\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  NnuM�����-z @@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@Ⅳ��@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@Ⅳ��ׁ��@M]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@Ù����@���@���@������@���  O�.Y�|��@k��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@Ù���Ƣ���@M������]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@ɕ��������@����������@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@ん�����@~@ɕ�ん�����M]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  P߆S!�'����@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@晉��@��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ȅ����M�����]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ׁ���M]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ׁ���㙅�M]^@@@@@@@@@@@@@@@@@@  Q�}������!��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉���م�M]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��㙁����M]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@�����@������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��  R��,����������������@@@@@@@Ó�����Ƣ���@M]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@\����@~@\��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  S�R�`������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@Ⅳ@ׁ��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���������  T7�V��U ��G�R����@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�Ⅳ��ׁ��@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�Ⅳ��ׁ��@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  U�}���v�3[@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@��@���������@~@}\����}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@����@�������@L~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���������@~@}\����������}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@  V�����9�ͱ@@@@@@@@����@�������@L~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���������@~@}\������������}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���������@~@}\������������}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  WH�D'��-w�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@����@���������@~@}\����������}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@  X��A��k����@ׁ��扄��@@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@ׁ��ȅ����@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@ז���≩�@@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@兙�◁��@@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@Ö��@@@@@@@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  Y}�zg�D��HT@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@Ӆ��ԁ����@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@㖗ԁ����@@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@����@���������@~@}\�����������}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@ׁ��扄��@@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@ׁ��ȅ  ZG�*%�Y�4ō����@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@ז���≩�@@~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@兙�◁��@@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@Ö��@@@@@@@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@Ӆ��ԁ����@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  [�n�*�m~���@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@㖗ԁ����@@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@����@���������@~@}\������������}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@ׁ��扄��@@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@ׁ��ȅ����@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@ז���≩�@@~@  \{:�2����U�4��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@兙�◁��@@~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@Ö��@@@@@@@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@Ӆ��ԁ����@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@㖗ԁ����@@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ]<a�w�Y�lض�s@@@@@@@@@@@@@@@@�������������@@@@@@@@@����@���������@~@}\������������}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@ׁ��扄��@@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@ׁ��ȅ����@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@ז���≩�@@~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@兙�◁��@@~@�^@@@@@  ^
w��D�4��h@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@Ö��@@@@@@@~@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@Ӆ��ԁ����@~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@㖗ԁ����@@~@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@����@���������@~@}\������}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  _h짂�!Q��@@@@@@@@@�������������@@@@@@@@@@@ׁ��扄��@@~@����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@ׁ��ȅ����@~@�����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@ז���≩�@@~@����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@兙�◁��@@~@����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@��@�Ö��@~@`�^@@@@@@@@@@@@@  `�����Ei�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@Ö��@~@�������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@Ö��@@@@@~@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  a���ҹМ�e@@�������������@@@@@@@@@@@Ӆ��ԁ����@~@�����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@㖗ԁ����@@~@����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@��@�֙����@~@}\���������}^@@@@@@@@@@@@  bM&u���W�܇@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@ׁ��扄��@@~@�ׁ��ȅ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@ׁ��ȅ����@~@�ׁ��扄��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�����  c`;�	~<��	X"��������@@@@@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�Ⅳ��ׁ��@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@Ù����@��@�����@���@������@����@@@@@@@@@@@@  d
G"�h�I��;J@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�Ù���Ƣ���@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�Ù���Ƣ���@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@������@@@@@@@@@@@@@@@@@@@@@@@����@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������������  e
�BTl�O=:$�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�Ɖ��Ձ��@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ř�Ԣ�@@@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  f����������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@Ɖ��Ձ��@~@l����M������]@N@�}��}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@È���@�������@������@����@������@��@���K@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@  g�"賩%��̠Y@��@~@����Ml����MƉ��Ձ��]@z@�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@Ɇ@⣙���@����@������k@����@������@���@������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@Ɇ@��@Ln@`�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@Ɇ@�����M��]@~@`�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  h'�Si�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@ř�Ԣ�@~@}�����M]@������K@}@N@����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@ŕ�Ɇ^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@Ɇ@������Ml����MƉ������]]@~@`�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@ř�Ԣ�@~@}������M]@������K@}@N@����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@ŕ��  i>��:�z�l��ִ�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@ŕ�Ɇ^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@��@������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@��@ř�Ԣ�@Ln@}@}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  j�A�M�;v�I<�@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@╄ׇ�Ԣ�@M}\������}z}Ù���Ƣ���}z@}@}@z@ř�Ԣ�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@ŕ���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@֗��MÙ����]@������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@��@~@����Ml��  k�����ЫŔ浄�MƉ������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@z@�m�����@N@�m������@N@�m�����@N@�m��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@z@�m�����@N@�m�����@z@���]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@Ɇ@��@~@`�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@ř�Ԣ�@~@}����M]@������K@}@N@����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  l�+��C�%C��q@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@ŕ�Ɇ^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@��@������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@��@ř�Ԣ�@Ln@}@}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@╄ׇ�Ԣ�@M}\�����  m�bk��[��O�}z}Ù���Ƣ���}z@}@}@z@ř�Ԣ�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@ŕ���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  n�4�jBӷB�C@@@@@@@@@@@@@�������������@@@@@�Ù���Ƣ���@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@晉��@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNN  o�FO]���GF�NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉��ā��@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉��ā��@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@¤����@@@@@@@@@@@@@@@@@@@@@@�����@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@Ӆ�@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  p���yg�z���@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@������@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@ħ�����@@@@@@@@@@@��@@@@@@@@@@@@@@@@@@�������M}m������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@\@  qy/]���%�@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�¨����@@@@@@@@@@@�@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ř�Ԣ�@@@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�  ro9�j�`ZmW�|������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@�������@��@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@������@Ml����M¤����]zl����Mん�����]zӅ�  s�z,2��»�eY]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@�����@����@��@������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@¨����@~@�����M��zl����M¤����]zӅ�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@Ɇ@¨����@Ln@Ӆ�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��������  t:�Y��������������@@@@@@@@@ř�Ԣ�@~@}�����M]@������K@}@N@����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@ŕ���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@��������@�����@��������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@�ֆ����@N~@¨����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  uR��fp)����c@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉��ā��@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@  v������2���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@晉��@������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉��ȅ����@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  wr���>l�/�C�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉��ȅ����@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@㉣��@@@@@@@@@@@@@@@@@@@@@@@@����@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@Ù������ā��@@@@�@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@œ  x��֮�M��H}҅����@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@�������@���@�������@���@����@ȉ�@�����@@@@@@@@@@@@@@@@@  y˵ �;�$� ���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}l���`�K�}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}l}@N@�}��������}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@��������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@Ӗ�������  z7y�@h�.�P�MtM�]@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}�@�@���}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}LL}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@Ù������ā��@~@l����Ml����M]z\����]Nl����Ml����M]z\����]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}aÙ������ā��@M�z}@N@Ù������ā��@N@}]}N@��z��]^@@@@@@@@@@  {-��f3M���@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}aי������@M�������@��K�@M����@���Ö���k@����]]}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@œ�����@~@}a㉣��@M}@N@l����M㉣��]@N@}]}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}nn}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}�����  |��F"˒ ��}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@����@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@Ӗ�������M�]@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}�@�@���}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  }9�w�1�[l۽�@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}LL}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}a㨗�@aÁ�����}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}aׁ���@�@�@�}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}nn}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}������}N��z�  ~�Ɇ5)����L]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@Ӗ�������M�]@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}�@�@���}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �E�ΐ���/�hG@@@@@@@@@@�������������@@@@@@@晉��ā��M}LL}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}a㨗�@aƖ��}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}a⤂����@a㨗��}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}aՁ��@a��}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@��@���������@~@}\���}^@@@@@@@@  ����16��Rf@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@Ɩ��@~@ą�����Ɩ��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@Ɩ��@~@���������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��LU#���Z�@@@�������������@@@@@@@œ�����@~@}a��Ɩ��@a}@N@l����MƖ��]@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}aŕ������@a払����ŕ������}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}nn}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}������}N��z�]^@@@@@@@@@@@@  �ޝ��q6q�g2@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@����@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@Ӗ�������M�]@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}�@�@���}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����  �c|j�i�ebY�����������@@@@@@@晉��ā��M}LL}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}@@aƖ��@LL@a��@�@�@�@nn}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}@@aי��Ⅳ@�@a���@aㅧ�@�}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}nn}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}������}N��z�]^@@@@@@@@@@@@@@@@@@@  �����w>w��Ȑ@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉��ȅ����@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�����������  �����G�I�eZ݀��@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@晉��@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉��ׁ���@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉��ׁ���@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �(qk@�G+�y��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@œ�����@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���⣙���@@@@@�@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@  �~����X8���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�@@@@@@@@@@@@@@@�@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�@@@@@@@@@@@@@@@�@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�@@@@@@@@@@@@@@@�@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@ׁ���������@@@@@�@@@@@@@@@@@@@@@@@@@}�M]}@@@@@@@@@@@@@@@@@  ��ZY ��FJG�H@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@ׄ�ㅧ�@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@����@  �)1Y���	�k����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@���@���@l���M��������]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@aa@����@�@���@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@�����������@~@⣁��ׁ��M]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ���z��x���Ò@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@aa@����@�@�����@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@����@��������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@���@���@l���M��������]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@晉��ā��M}M}z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@ׄ�ㅧ�@  ����jrj�p&�T~@����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@aa@������@�����������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@���@�@~@�@��@l���Mׁ���������]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@�@~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@�@~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �1��F?�fip�@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@���@�@~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@�@~@l����Ml�����Mׁ���������z�z�]zl�����Mׄ�ㅧ�z�N�]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@��@�@n@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@�@N~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@ׄ�ㅧ�@~  ��e�6b%��M�,@l�������M}�}zׄ�ㅧ�z�z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@�@N~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �8g�j�RPGtR@@@@@@@@@@@@@@�������������@@@@@@@@@@@aa@�����@�����@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@晉��ā��Ml�����Mׄ�ㅧ�]zl���Ml�����Mׄ�ㅧ�]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@晉��ā��M}]}}}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@aa@����@����@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@����@��������^@@@@@@@@  �o�fBϦ�[b��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@��@���@l���M��������]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@aa@������@����@�����������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@����@����@~@}�}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �n�9��+��b�@@@@@@@�������������@@@@@@@@@@@@@@@@@ŕ�ׁ��M�����������]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@�����������@~@⣁��ׁ��M]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@����@����@~@}�}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@晉��ā��M}M]}}}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@����@����@~@}`}^@@@@@@@@@  �����%]�{@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@晉��ā��M}M]}}}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@晉��ā��M}M]}}}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ���N�q����>B��������������@@@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@aa@�����@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@ŕ�ׁ��M�����������]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��j([�L�;Sk@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@�����@��������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉��ׁ���@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������  �ubۚ�SA<������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@⣁��@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�⣁��ׁ��@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��+�so_F����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�⣁��ׁ��@@@@@@@@��@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@����ז�@@@@@@@@@�@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@œ�����@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@  �
I���,�9�2_�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@�ւ����@N~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��+��w��J��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@Ӗ�������M�ւ����]@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@����Ֆ@N~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@ׁ��ւ����M����Ֆ]@~@�ւ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@œ�����@~@l����M�ւ����]@N@}@�@���}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@�  �ʢO���^���♉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}LL}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}a㨗�@aׁ��}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}aׁ����@�@�@�}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}aم�������@�@�@�}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@  ��B�}y�E@|j@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@�ւ����@N~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@œ�����@~@}aÖ������@}@N@l����M�ւ����]@N@}@�@�}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}nn}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā�  ����ڥ���O��M}������}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@Ӗ�������M�ւ����]@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@œ�����@~@l����M�ւ����]@N@}@�@���}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@  ���wE-�P��@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}LL}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@œ�����@~@}aӅ����@}@N@l����M�ւ����@N@�]@N@}@�@�}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@  ��aĸ�gB�	�C�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}nn}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}������}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@����ז�@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �o�#� d��H��@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@��@�����@�@����@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}��}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@���@�������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@œ�����@~@}a��@}@N@l��  ����%��-�2���M�����≩�]@N@}@�}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@���@�������@M�k�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@œ�����@~@}�@�@�@�@}@N@l����M����ԁ����]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �HD�;��3�I��@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@}@}@N@l����M����ȅ����@`@���ԁ����]@N@}@�}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@���@��������@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@œ�����@~@l����M����◁��]@N@  ���ӱ�c�e`���}@��}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@������@����ז�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �ܸ������ld�@@@@�������������@@@@@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�⣁��ׁ��@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@ŕ�@����@@@@@@@@@@@@@@@@@@@@@@@@@@  �X&���sB�{ɣ@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ŕ�ׁ��@@@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ŕ�ׁ��@@@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@⣙���⣁��@@@@@@@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���  �%؆�w�Y�bHL�����������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@œ�����@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@⣙���ŕ�@@@@@@@�@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �ș,P9��KR��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@aa@��@����@���@����@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@晉��ā��M}��}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@������ŕ�@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@晉��ā��M}���������}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@����������  ��P_2N��b�����@@@@@@@@@晉��ā��M}������}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@�ւ����@N~@�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@Ӗ�������M�ւ����]@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �,�X��w�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@œ�����@~@l����M�ւ����]@N@}@�@���}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@œ�����@~@l����M⣙���ŕ�@`@������⣁��]@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@  �h)��%��8�4@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@晉��ā��M}������}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �f�
D�T��&�� @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ŕ�ׁ��@@@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@晉��@�����@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNN  �`Մ�[�Ug�l��NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉��ׁ���㙅�@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉��ׁ���㙅�@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�@@@@@@@@@@@@@@@�@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �Cv|������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@œ�����@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@  �CI�������.�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@Ӗ�������M�]@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}�@�@���}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}LL}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}a㨗�@aׁ���}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �JU�گ�0��˼@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@������@����@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@œ�����@~@}aÖ���@}@N@l����M����Ֆ]@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@  ��3���/hL�
b@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@������@���������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@œ�����@~@}aԅ����@�@�@�@}@N@l����M����扄��]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@}@}@N@l����M����ȅ����]@N@}@�}@N��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �7	P���vi`{�C@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@������@������@���������@��@����@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}a҉��@�}z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@���@�@~@�@��@����Ֆ^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@��@l���M�z��]@~@�^@@@@@  �i̙��fF��6�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@晉��ā��M��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@œ�����@~@}@}@N@l����Mׁ��ւ����M�]]@N@}@�@�}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��hX����d�4��@@@@@@@@�������������@@@@@@@������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}@�}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}nn}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}������}N��z�]^@@@@@@@  �W7��i��~��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉��ׁ���㙅�@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ���Vn!���:D@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@晉��@�م�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉���م�@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉���م�@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@  �.��A�wC��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�@@@@@@@@@@@@@@@�@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@œ�����@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������  ��%|]���Z�������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@�����@�م�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@�م�@~@�ֆ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �6���:t:�s�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}����}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@KKK@������@��@�������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@œ�����@~@}�@}@N@l����M�ւ����@N@�]@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������  ����D���!�@@@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@KKK@����@�����@`@����@��@������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@œ�����@~@}����������@�����@�@}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@  ��@(��"�t<E�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@KKK@�م�@�������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@���@�@~@�@��@�ւ����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@œ�����@~@l����Ml�����Ml���MӖ�������M�]z��z�]z}�}]]@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@  ����H*�H�.�@@@@@@@@@@@}@�����@�@}@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��*���df��z�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉���م�@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@晉��@�������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNN  ��b�;�'K6�\�hNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉��㙁����@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉��㙁����@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@œ�����@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ���@�m�%�n��@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}�������}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}LL}  ��1�P$�J��9N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@�����@������@��@�������@��@�م�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@œ�����@~@}a≩�@}@N@l����M�ւ����@N@�]@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��:��Q��B�%�@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}aٖ��@�@�@�}N��z��]^@@@@@aa@���������@��@Á�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}aɕ��@�@�@�}N��z��]^@@@@@aa@���������@��@ɕ��@����������@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}nn}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@aa@������@��@�م�@@@@  �sp=3B`~쁀�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}���������}N��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@œ�����@~@l����M�م�]@N@��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��Mœ�����zl���Ml�����Mœ�����]]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �z�80�5�yKĲ�@@@@@@@@@@@@�������������@@@@@@@aa@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@晉��ā��M}ll���}N��z�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�晉��㙁����@@@@@�@@@@@@@@@@@  � #��?!���8g�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@Ó���@���@������@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@  �wz[�U��}`�8@@@@@�������������@@@@@�Ó�����Ƣ���@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�Ó�����Ƣ���@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ř�Ԣ�@@@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �o
+<�z9��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@Ɇ@�����M��]@~@`�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@ř�Ԣ�@~@}�����M]@������K@}@N@����������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@╄ׇ�Ԣ�@M}\������}z}Ó���Ƣ���}z@}@}@z@ř�Ԣ�]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@ŕ�Ɇ^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@��  �x�1zd����P�����������@@@@@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�Ó�����Ƣ���@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN  ĩ��l���RNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@ɕ��������@あ��@ł����@`n@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ɕ�ん�����@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ɕ�ん�����@@@@@@��@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@���������  ����w�R��%�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@Ö�����@�@Ǚ�����@È�������@⣙���@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@��������@@@@@@@@@@��@@@@@@@@@@@@@@@@@@������M}�������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@������@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@  �nuW8�@
�~�V@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@��@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@������@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@  Ǒ`�ى
s���b@@�@������@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@��@@@@@@@@@@@@@@@@@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@  �cZ��j)(�[KL@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@���������@@@@@@@@@��@@@@@@@@@@@@@@@@@@������M}��������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@��������@@@@@@@@@@@@@@@@@@@@����@@@@�������M\�������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���  �%{r�Fg���"�r�¨���@@@@@@@@@@@@@@@@@@@@@@��@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@����Ɩ����@@@@@@@@@@@@@@@@@@@@��@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@����і�Ձ��@@@@@@@@@@@@@@@@@@@��@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@����і�ɕ�@@@@@@@@@@@@@@@@@@@@��@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���ř���@@@@@@@@@@@@@@@@@@@@@���@@@@�������M\�������]@@@@@@@@@@  �3��FB�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@��������@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@�����@@@@@@@@@@@@@@@@@@@@@@@@@��@�@�������M��������z���]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@����������@������@���@�������@���@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�ん�����@@@  ˔�̍WqAT�d�5@@@@@@�@@@@@@@@@@@@���@@@@���M\����}��}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�んł����@@@@@@@@�@@@@@@@@@@@@���@@@@���M\����}��}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@���@@@@@@@@@@@@@@@�@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@���@@@@@@@@@@@@@@@�@@@@@@@@@@@@@���@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@���@@@@@@@@@@@@@@@�@@@@@@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �i��]�����E@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@����������@������@`@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@��偓��@@@@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@�偓��@@@@@@@@@@@@@@@@@@@@@@@@@��@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@  ͪ�&Mk�&��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@aa@���@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@��������@M��������zl���M��������]z}��������}z}\}z}@}z�����]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@aa@������@�@����������@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ΀"��*t�R�v@@@@@@@@@@@@@@@@�������������@@@@@@@@���@�偓��@~@�@��@���^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@l�����Mんł����z�偓��N�z�]@~@�偓��^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@aa@������@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@�������@M�����z�zんł�  ��)�M(4���b���z���z���z�z�z���zん�����z��z��z��]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@aa@������@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@������@ん�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��֞c���`��(�@@@@@@@@@�������������@@@@@�ɕ�ん�����@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@ǅ�@�@�����@����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN  ш�m+�Os�#�[NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@ׇ���������@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@ć���������@@@@@@@��@@@@@@@@@@@���@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@ć�������@@@@@@@@@��@@@@@@@@@@@@@@\@@@�������M}mm�����}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@Ģ�������@@@@@@@@@��@@@@@@@@@@@@@@\@@@�������M}��������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ҮP)*x���B9@@�������������@@@@@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@���@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@ą�����@@@@@@@@@@@�@@@@@@@@@@@@@���@�@�����M������m�]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@������m�@~@��������^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@م����@l����Ml�����M������@z@}�}]]@N@}  Ӏ c�ך=L�%@z@}@N@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@l���M��������M������]]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@ׇ���������@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�����  �W�F�J�<�Wem��������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aa@⅕�@י�����@ԅ�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@aaNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�╄ׇ�Ԣ�@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�╄ׇ�Ԣ�@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@  ��,7	�h�]X�?W@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���㨗�@@@@@@@@@@@@@@@@@@@@@@@���@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@��������@@@@@@@@@@@@@@@@@@@@@@���@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���Ʉ@@@@@@@@@@@@@@@@@@@@@@@@@@��@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���ř�@@@@@@@@@@@@@@@@@@@@@@@����@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@������������  ։��P�K�ϬD�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@��������@@@@@@@@��@@@@@@@@@@@@@@@@@@������M}��������}]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@ԅ�����Ʉ@@@@@@@@@@@@@@@@@@@@@�@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@ԅ�����Ɖ��@@@@@@@@@@@@@@@@@@��@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@ԅ�����ā��@@@@@@@@@@@@@@@@@���@@@@�����@�������M\�  �qK��9�9 �%(
������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@ԅ�����ā���@@@@@@@@@@@@@@@@@@��@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@ԅ�����㨗�@@@@@@@@@@@@@@@@@@��@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@Á��⣒ŕ���@@@@@@@@@@@@@@@@���@@@@�����@�������M\�������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@Á��⣒Ö���@@@@@@@@@@@@@@@@@@��@�@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�  �؈�����|7
�R@@ԅ�����҅�@@@@@@@@@@@@@@@@@@@@�@@@@�����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@@���ř���@@@@@@@@@@@@@@@@@@@@���@@@@�������M\�������]@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@��Ԣ�@@@@@@@@@@@�@@@@@@@@@@@@@@��@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�@���Ԣ�@@@@@@@@@@�@@@@@@@@@@@@����@@@@@@@@@@@@@@@@@@@@@@@@@@  ����9+��h@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@��@���Ʉ@Ln@}@}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@��Ԣ  �0���y�6UF�D�@@~@���Ʉ^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@���Ԣ�@~@���ř�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@��@���㨗�@~@}\������}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@��Ԣ�@@~@}�������}^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  �T�X�+�S�p@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@���Ԣ�@~@}ř���@}@N@l�����M��������]@N@}@z@}@N@���ř�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@���Ԣ�@~@���ř�^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@�����^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@�����^@@@@@@@  ��aG���x�e�Jw@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@��������@M��Ԣ�z@}�������@@@����}@z@���Ԣ�@z@l���M���Ԣ�]@z@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@���㨗�@z@}\������}@z@�@z@}@}@z@�����]^@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ݳ.�$l����@@@@@@@@@@@@@@@@@@@@�������������@@@@@@a���`����@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@�������������@@@@@�╄ׇ�Ԣ�@@@@@@@@�@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                                                                                                                                                                                                                                                                            �����u�Ay�>                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ߉s�Xo  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ����x�I�x����[  ���:%�hQk �